-- code generated from the following source code:
--   stdlib.ecl
--   ../benchs/queens/nqueens.ecl
--
-- with the following command:
--
--    ./eclat ../benchs/queens/nqueens.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal argument : in value(0 to 11);
       signal result : out value(0 to 57));
       
end entity;
architecture rtl of main is

  type t_state is (IDLE405);
  signal \state%now\, \state%next\: t_state;
  type t_state_var609 is (IDLE444, PAUSE_SET445, Q_WAIT446);
  signal \state_var609%now\, \state_var609%next\: t_state_var609;
  type t_state_var608 is (IDLE450, PAUSE_GET451, Q_WAIT452);
  signal \state_var608%now\, \state_var608%next\: t_state_var608;
  type t_state_var607 is (IDLE420, \$1594\, \$1607_LOOP99401\, \$1619_LOOP99398\, \$1633_LOOP99399\, \$1646_LOOP99400\, PAR454, PAUSE_GET457, PAUSE_SET421, Q_WAIT422, Q_WAIT458);
  signal \state_var607%now\, \state_var607%next\: t_state_var607;
  type t_state_var606 is (IDLE486, PAUSE_SET487, Q_WAIT488);
  signal \state_var606%now\, \state_var606%next\: t_state_var606;
  type t_state_var605 is (IDLE492, PAUSE_GET493, Q_WAIT494);
  signal \state_var605%now\, \state_var605%next\: t_state_var605;
  type t_state_var604 is (IDLE462, \$1660\, \$1673_LOOP99401\, \$1685_LOOP99398\, \$1699_LOOP99399\, \$1712_LOOP99400\, PAR496, PAUSE_GET499, PAUSE_SET463, Q_WAIT464, Q_WAIT500);
  signal \state_var604%now\, \state_var604%next\: t_state_var604;
  type t_state_var603 is (IDLE528, PAUSE_SET529, Q_WAIT530);
  signal \state_var603%now\, \state_var603%next\: t_state_var603;
  type t_state_var602 is (IDLE534, PAUSE_GET535, Q_WAIT536);
  signal \state_var602%now\, \state_var602%next\: t_state_var602;
  type t_state_var601 is (IDLE504, \$1726\, \$1739_LOOP99401\, \$1751_LOOP99398\, \$1765_LOOP99399\, \$1778_LOOP99400\, PAR538, PAUSE_GET541, PAUSE_SET505, Q_WAIT506, Q_WAIT542);
  signal \state_var601%now\, \state_var601%next\: t_state_var601;
  type t_state_var600 is (IDLE570, PAUSE_SET571, Q_WAIT572);
  signal \state_var600%now\, \state_var600%next\: t_state_var600;
  type t_state_var599 is (IDLE576, PAUSE_GET577, Q_WAIT578);
  signal \state_var599%now\, \state_var599%next\: t_state_var599;
  type t_state_var598 is (IDLE546, \$1792\, \$1805_LOOP99401\, \$1817_LOOP99398\, \$1831_LOOP99399\, \$1844_LOOP99400\, PAR580, PAUSE_GET583, PAUSE_SET547, Q_WAIT548, Q_WAIT584);
  signal \state_var598%now\, \state_var598%next\: t_state_var598;
  type t_state_var597 is (IDLE409, \$1588\, \$1857\, PAR586, PAUSE_GET410, PAUSE_SET588, PAUSE_SET591, Q_WAIT411, Q_WAIT589, Q_WAIT592);
  signal \state_var597%now\, \state_var597%next\: t_state_var597;
  type array_value_32 is array (natural range <>) of value(0 to 31);
  signal \$1209_src\ : array_value_32(0 to 7);
  signal \$$1209_src_value\ : value(0 to 31) := (others => '0');
  signal \$$1209_src_ptr\ : natural range 0 to 7 := 0;
  signal \$$1209_src_ptr_write\ : natural range 0 to 7 := 0;
  signal \$$1209_src_write\ : value(0 to 31) := (others => '0');
  signal \$$1209_src_write_request\ : std_logic := '0';
  signal \$1216_dst\ : array_value_32(0 to 7);
  signal \$$1216_dst_value\ : value(0 to 31) := (others => '0');
  signal \$$1216_dst_ptr\ : natural range 0 to 7 := 0;
  signal \$$1216_dst_ptr_write\ : natural range 0 to 7 := 0;
  signal \$$1216_dst_write\ : value(0 to 31) := (others => '0');
  signal \$$1216_dst_write_request\ : std_logic := '0';
  signal \$1217_r\ : array_value_32(0 to 0);
  signal \$$1217_r_value\ : value(0 to 31) := (others => '0');
  signal \$$1217_r_ptr\ : natural range 0 to 0 := 0;
  signal \$$1217_r_ptr_write\ : natural range 0 to 0 := 0;
  signal \$$1217_r_write\ : value(0 to 31) := (others => '0');
  signal \$$1217_r_write_request\ : std_logic := '0';
  signal \$1614%next\, \$1614%now\, \$1812%next\, \$1812%now\, \$1690%next\, 
         \$1690%now\, \$1704%next\, \$1704%now\, \$1709%next\, \$1709%now\, 
         \$1770%next\, \$1770%now\, \$1706%next\, \$1706%now\, \$1717%next\, 
         \$1717%now\, \$1615%next\, \$1615%now\, \$1810%next\, \$1810%now\, 
         \$1636%next\, \$1636%now\, \$1655%next\, \$1655%now\, \$1808%next\, 
         \$1808%now\, \$1616%next\, \$1616%now\, \$1784%next\, \$1784%now\, 
         \$1758%next\, \$1758%now\, \$1722%next\, \$1722%now\, \$1838%next\, 
         \$1838%now\, \$1836%next\, \$1836%now\, \$1820%next\, \$1820%now\, 
         \$1772%next\, \$1772%now\, \$1746%next\, \$1746%now\, \$1680%next\, 
         \$1680%now\, \$1721%next\, \$1721%now\, \$1813%next\, \$1813%now\, 
         \$1760%next\, \$1760%now\, \$1656%next\, \$1656%now\, \$1643%next\, 
         \$1643%now\, \$1759%next\, \$1759%now\, \$1754%next\, \$1754%now\, 
         \$1610%next\, \$1610%now\, \$1857_arg%next\, \$1857_arg%now\, 
         \$1769%next\, \$1769%now\, \$1641%next\, \$1641%now\, \$1786%next\, 
         \$1786%now\, \$1654%next\, \$1654%now\, \$1822%next\, \$1822%now\, 
         \$1688%next\, \$1688%now\, \$1773%next\, \$1773%now\, \$1785%next\, 
         \$1785%now\, \$1612%next\, \$1612%now\, \$1774%next\, \$1774%now\, 
         \$1749%next\, \$1749%now\, \$1720%next\, \$1720%now\, \$1757%next\, 
         \$1757%now\, \$1652%next\, \$1652%now\, \$1651%next\, \$1651%now\, 
         \$1839%next\, \$1839%now\, \$1624%next\, \$1624%now\, \$1650%next\, 
         \$1650%now\, \$1747%next\, \$1747%now\, \$1695%next\, \$1695%now\, 
         \$1824%next\, \$1824%now\, \$1626%next\, \$1626%now\, \$1823%next\, 
         \$1823%now\, \$1748%next\, \$1748%now\, \$1708%next\, \$1708%now\, 
         \$1761%next\, \$1761%now\, \$1826%next\, \$1826%now\, \$1849%next\, 
         \$1849%now\, \$1809%next\, \$1809%now\, \$1783%next\, \$1783%now\, 
         \$1679%next\, \$1679%now\, \$1847%next\, \$1847%now\, \$1689%next\, 
         \$1689%now\, \$1642%next\, \$1642%now\, \$1796%next\, \$1796%now\, 
         \$1718%next\, \$1718%now\, \$1598%next\, \$1598%now\, \$1768%next\, 
         \$1768%now\, \$1841%next\, \$1841%now\, \$1629%next\, \$1629%now\, 
         \$1775%next\, \$1775%now\, \$1840%next\, \$1840%now\, \$1694%next\, 
         \$1694%now\, \$1781%next\, \$1781%now\, \$1854%next\, \$1854%now\, 
         \$1788%next\, \$1788%now\, \$1743%next\, \$1743%now\, \$1851%next\, 
         \$1851%now\, \$1617%next\, \$1617%now\, \$1827%next\, \$1827%now\, 
         \$1715%next\, \$1715%now\, \$1837%next\, \$1837%now\, \$1653%next\, 
         \$1653%now\, \$1676%next\, \$1676%now\, \$1692%next\, \$1692%now\, 
         \$1742%next\, \$1742%now\, \$1848%next\, \$1848%now\, \$1745%next\, 
         \$1745%now\, \$1625%next\, \$1625%now\, \$1702%next\, \$1702%now\, 
         \$1716%next\, \$1716%now\, \$1691%next\, \$1691%now\, \$1693%next\, 
         \$1693%now\, \$1835%next\, \$1835%now\, \$1611%next\, \$1611%now\, 
         \$1622%next\, \$1622%now\, \$1825%next\, \$1825%now\, \$1623%next\, 
         \$1623%now\, \$1649%next\, \$1649%now\, \$1782%next\, \$1782%now\, 
         \$1681%next\, \$1681%now\, \$1850%next\, \$1850%now\, \$1678%next\, 
         \$1678%now\, \$1853%next\, \$1853%now\, \$1705%next\, \$1705%now\, 
         \$1787%next\, \$1787%now\, \$1852%next\, \$1852%now\, \$1639%next\, 
         \$1639%now\, \$1628%next\, \$1628%now\, \$1771%next\, \$1771%now\, 
         \$1815%next\, \$1815%now\, \$1638%next\, \$1638%now\, \$1677%next\, 
         \$1677%now\, \$1755%next\, \$1755%now\, \$1814%next\, \$1814%now\, 
         \$1707%next\, \$1707%now\, \$1578%next\, \$1578%now\, \$1613%next\, 
         \$1613%now\, \$1627%next\, \$1627%now\, \$1640%next\, \$1640%now\, 
         \$1821%next\, \$1821%now\, \$1703%next\, \$1703%now\, \$1811%next\, 
         \$1811%now\, \$1719%next\, \$1719%now\, \$1756%next\, \$1756%now\, 
         \$1730%next\, \$1730%now\, \$1637%next\, \$1637%now\, \$1683%next\, 
         \$1683%now\, \$1834%next\, \$1834%now\, \$1682%next\, \$1682%now\, 
         \$1744%next\, \$1744%now\, \$1664%next\, \$1664%now\ : value(0 to 32) := (others => '0');
  signal \$1594_arg%next\, \$1594_arg%now\, \$1726_arg%next\, 
         \$1726_arg%now\, \$1660_arg%next\, \$1660_arg%now\, 
         \$1792_arg%next\, \$1792_arg%now\, \$1592%next\, \$1592%now\ : value(0 to 3) := (others => '0');
  signal \result403%next\, \result403%now\ : value(0 to 57) := (others => '0');
  signal \$1751_loop99398_id%next\, \$1751_loop99398_id%now\, 
         \$1831_loop99399_id%next\, \$1831_loop99399_id%now\, 
         \$1633_loop99399_id%next\, \$1633_loop99399_id%now\, 
         \$1805_loop99401_id%next\, \$1805_loop99401_id%now\, 
         \$1699_loop99399_id%next\, \$1699_loop99399_id%now\, 
         \$1619_loop99398_id%next\, \$1619_loop99398_id%now\, 
         \$1844_loop99400_id%next\, \$1844_loop99400_id%now\, 
         \$1588_id%next\, \$1588_id%now\, \$1778_loop99400_id%next\, 
         \$1778_loop99400_id%now\, \$1607_loop99401_id%next\, 
         \$1607_loop99401_id%now\, \$1739_loop99401_id%next\, 
         \$1739_loop99401_id%now\, \$1685_loop99398_id%next\, 
         \$1685_loop99398_id%now\, \$1857_id%next\, \$1857_id%now\, 
         \$1673_loop99401_id%next\, \$1673_loop99401_id%now\, 
         \$1792_id%next\, \$1792_id%now\, \$1726_id%next\, \$1726_id%now\, 
         \$1594_id%next\, \$1594_id%now\, \$1817_loop99398_id%next\, 
         \$1817_loop99398_id%now\, \$1660_id%next\, \$1660_id%now\, 
         \$1712_loop99400_id%next\, \$1712_loop99400_id%now\, 
         \$1765_loop99399_id%next\, \$1765_loop99399_id%now\, 
         \$1646_loop99400_id%next\, \$1646_loop99400_id%now\ : value(0 to 11) := (others => '0');
  signal \$1588_arg%next\, \$1588_arg%now\ : value(0 to 64) := (others => '0');
  signal \$1861%next\, \$1861%now\, \$1577_o%next\, \$1577_o%now\ : value(0 to 127) := (others => '0');
  signal \$$1217_r_lock%next\, \$$1217_r_lock%now\, \$$1216_dst_lock%next\, 
         \$$1216_dst_lock%now\, \$$1209_src_lock%next\, 
         \$$1209_src_lock%now\, \$v412%next\, \$v412%now\, \rdy503%next\, 
         \rdy503%now\, \$1600%next\, \$1600%now\, \$1606%next\, \$1606%now\, 
         \$v518%next\, \$v518%now\, \$v510%next\, \$v510%now\, \$v474%next\, 
         \$v474%now\, \$1799%next\, \$1799%now\, \$1711%next\, \$1711%now\, 
         \$v523%next\, \$v523%now\, \rdy533%next\, \rdy533%now\, 
         \$v594%next\, \$v594%now\, \$1763%next\, \$1763%now\, \$v519%next\, 
         \$v519%now\, \$1658%next\, \$1658%now\, \$1579%next\, \$1579%now\, 
         \$1738%next\, \$1738%now\, \$v558%next\, \$v558%now\, \$1764%next\, 
         \$1764%now\, \$v556%next\, \$v556%now\, \$1660_result%next\, 
         \$1660_result%now\, \$1801%next\, \$1801%now\, \rdy575%next\, 
         \rdy575%now\, \$v468%next\, \$v468%now\, \$1605%next\, \$1605%now\, 
         \$v587%next\, \$v587%now\, \$1580_led%next\, \$1580_led%now\, 
         \$v455%next\, \$v455%now\, \$v514%next\, \$v514%now\, \$v582%next\, 
         \$v582%now\, \$1631%next\, \$1631%now\, \$v477%next\, \$v477%now\, 
         \$v475%next\, \$v475%now\, \rdy443%next\, \rdy443%now\, 
         \$v560%next\, \$v560%now\, \result526%next\, \result526%now\, 
         \$1668%next\, \$1668%now\, \$v522%next\, \$v522%now\, \$1586%next\, 
         \$1586%now\, \$v437%next\, \$v437%now\, \$v564%next\, \$v564%now\, 
         \$v508%next\, \$v508%now\, \$v531%next\, \$v531%now\, \$v465%next\, 
         \$v465%now\, \$1804%next\, \$1804%now\, \rdy449%next\, \rdy449%now\, 
         \$1857_result%next\, \$1857_result%now\, \$1798%next\, \$1798%now\, 
         \rdy545%next\, \rdy545%now\, \$v430%next\, \$v430%now\, 
         \$1582%next\, \$1582%now\, \$v551%next\, \$v551%now\, \$v439%next\, 
         \$v439%now\, \$v515%next\, \$v515%now\, \$1733%next\, \$1733%now\, 
         \$1829%next\, \$1829%now\, \$v423%next\, \$v423%now\, \$v585%next\, 
         \$v585%now\, \$v549%next\, \$v549%now\, \$v563%next\, \$v563%now\, 
         \$v453%next\, \$v453%now\, \$1671%next\, \$1671%now\, \$1777%next\, 
         \$1777%now\, \$1667%next\, \$1667%now\, \$v498%next\, \$v498%now\, 
         \$v552%next\, \$v552%now\, \$1726_result%next\, \$1726_result%now\, 
         \$v554%next\, \$v554%now\, \$1800%next\, \$1800%now\, \$v479%next\, 
         \$v479%now\, \$1602%next\, \$1602%now\, \$v434%next\, \$v434%now\, 
         \$v472%next\, \$v472%now\, \$v436%next\, \$v436%now\, \$v489%next\, 
         \$v489%now\, \$v537%next\, \$v537%now\, \result442%next\, 
         \result442%now\, \$v397%next\, \$v397%now\, \$v426%next\, 
         \$v426%now\, \$v456%next\, \$v456%now\, \$1584%next\, \$1584%now\, 
         \$v424%next\, \$v424%now\, \$v555%next\, \$v555%now\, \$v438%next\, 
         \$v438%now\, \$v476%next\, \$v476%now\, \$v521%next\, \$v521%now\, 
         \$1632%next\, \$1632%now\, \$1792_result%next\, \$1792_result%now\, 
         \$v459%next\, \$v459%now\, \rdy485%next\, \rdy485%now\, 
         \$v509%next\, \$v509%now\, \rdy527%next\, \rdy527%now\, 
         \$v480%next\, \$v480%now\, \$v429%next\, \$v429%now\, \rdy404%next\, 
         \rdy404%now\, \rdy461%next\, \rdy461%now\, \$v565%next\, 
         \$v565%now\, \$v520%next\, \$v520%now\, \rdy419%next\, \rdy419%now\, 
         \$v573%next\, \$v573%now\, \$v435%next\, \$v435%now\, \$v593%next\, 
         \$v593%now\, \$v501%next\, \$v501%now\, \$v562%next\, \$v562%now\, 
         \$v466%next\, \$v466%now\, \$v467%next\, \$v467%now\, \$v473%next\, 
         \$v473%now\, \$v428%next\, \$v428%now\, \$v516%next\, \$v516%now\, 
         \$1587%next\, \$1587%now\, \$v478%next\, \$v478%now\, \$v590%next\, 
         \$v590%now\, \$1581%next\, \$1581%now\, \result418%next\, 
         \result418%now\, \$1830%next\, \$1830%now\, \$v432%next\, 
         \$v432%now\, \$1601%next\, \$1601%now\, \$v481%next\, \$v481%now\, 
         \$v495%next\, \$v495%now\, \$v433%next\, \$v433%now\, \$v559%next\, 
         \$v559%now\, \$v431%next\, \$v431%now\, \$v395%next\, \$v395%now\, 
         \$1669%next\, \$1669%now\, \$v470%next\, \$v470%now\, \$v469%next\, 
         \$v469%now\, \$1724%next\, \$1724%now\, \$1734%next\, \$1734%now\, 
         \$1583%next\, \$1583%now\, \$v497%next\, \$v497%now\, \$v539%next\, 
         \$v539%now\, \$1856%next\, \$1856%now\, \$1790%next\, \$1790%now\, 
         \$1672%next\, \$1672%now\, \result568%next\, \result568%now\, 
         \$1603%next\, \$1603%now\, \$v425%next\, \$v425%now\, 
         \$1594_result%next\, \$1594_result%now\, \$1697%next\, \$1697%now\, 
         \$v471%next\, \$v471%now\, \$1585%next\, \$1585%now\, \$1732%next\, 
         \$1732%now\, \$v427%next\, \$v427%now\, \$v581%next\, \$v581%now\, 
         \$1860%next\, \$1860%now\, \rdy408%next\, \rdy408%now\, 
         \rdy491%next\, \rdy491%now\, \$v543%next\, \$v543%now\, 
         \$v517%next\, \$v517%now\, \$v540%next\, \$v540%now\, \$v513%next\, 
         \$v513%now\, \result484%next\, \result484%now\, \$1843%next\, 
         \$1843%now\, \$v406%next\, \$v406%now\, \$v507%next\, \$v507%now\, 
         \result544%next\, \result544%now\, \$v550%next\, \$v550%now\, 
         \result502%next\, \result502%now\, \$v512%next\, \$v512%now\, 
         \result460%next\, \result460%now\, \$1645%next\, \$1645%now\, 
         \$v553%next\, \$v553%now\, \$v413%next\, \$v413%now\, \$v557%next\, 
         \$v557%now\, \$v579%next\, \$v579%now\, \$v561%next\, \$v561%now\, 
         \$1735%next\, \$1735%now\, \$1698%next\, \$1698%now\, \$1803%next\, 
         \$1803%now\, \$1666%next\, \$1666%now\, \$v447%next\, \$v447%now\, 
         \$v596%next\, \$v596%now\, \$v511%next\, \$v511%now\, \$1737%next\, 
         \$1737%now\, \rdy569%next\, \rdy569%now\ : value(0 to 0) := (others => '0');
  signal \$1619_loop99398_result%next\, \$1619_loop99398_result%now\, 
         \$1789_nb2%next\, \$1789_nb2%now\, \$1731_n%next\, \$1731_n%now\, 
         \$1663_i%next\, \$1663_i%now\, \$1604%next\, \$1604%now\, 
         \$1765_loop99399_result%next\, \$1765_loop99399_result%now\, 
         \result532%next\, \result532%now\, \$1795_i%next\, \$1795_i%now\, 
         \$1618_nb2%next\, \$1618_nb2%now\, \$1729_i%next\, \$1729_i%now\, 
         \$1805_loop99401_result%next\, \$1805_loop99401_result%now\, 
         \$1630_nb2%next\, \$1630_nb2%now\, \$1588_result%next\, 
         \$1588_result%now\, \result490%next\, \result490%now\, 
         \$1828_nb2%next\, \$1828_nb2%now\, \$1723_nb2%next\, 
         \$1723_nb2%now\, \$1842_nb2%next\, \$1842_nb2%now\, 
         \$1699_loop99399_result%next\, \$1699_loop99399_result%now\, 
         \$1802%next\, \$1802%now\, \$1646_loop99400_result%next\, 
         \$1646_loop99400_result%now\, \$1673_loop99401_result%next\, 
         \$1673_loop99401_result%now\, \$1739_loop99401_result%next\, 
         \$1739_loop99401_result%now\, \$1599_n%next\, \$1599_n%now\, 
         \$1778_loop99400_result%next\, \$1778_loop99400_result%now\, 
         \result407%next\, \result407%now\, \$1607_loop99401_result%next\, 
         \$1607_loop99401_result%now\, \$1844_loop99400_result%next\, 
         \$1844_loop99400_result%now\, \$1817_loop99398_result%next\, 
         \$1817_loop99398_result%now\, \$1855_nb2%next\, \$1855_nb2%now\, 
         \$1696_nb2%next\, \$1696_nb2%now\, \$1644_nb2%next\, 
         \$1644_nb2%now\, \$1657_nb2%next\, \$1657_nb2%now\, 
         \$1712_loop99400_result%next\, \$1712_loop99400_result%now\, 
         \result448%next\, \result448%now\, \$1750_nb2%next\, 
         \$1750_nb2%now\, \$1659_i%next\, \$1659_i%now\, \$1670%next\, 
         \$1670%now\, \$1776_nb2%next\, \$1776_nb2%now\, \$1591_x%next\, 
         \$1591_x%now\, \$1751_loop99398_result%next\, 
         \$1751_loop99398_result%now\, \$1725_i%next\, \$1725_i%now\, 
         \$1736%next\, \$1736%now\, \$1710_nb2%next\, \$1710_nb2%now\, 
         \$1831_loop99399_result%next\, \$1831_loop99399_result%now\, 
         \$1593_i%next\, \$1593_i%now\, \$1597_i%next\, \$1597_i%now\, 
         \$1665_n%next\, \$1665_n%now\, \$1791_i%next\, \$1791_i%now\, 
         \$1816_nb2%next\, \$1816_nb2%now\, \$1684_nb2%next\, 
         \$1684_nb2%now\, \result574%next\, \result574%now\, 
         \$1685_loop99398_result%next\, \$1685_loop99398_result%now\, 
         \$1797_n%next\, \$1797_n%now\, \$1633_loop99399_result%next\, 
         \$1633_loop99399_result%now\, \$1762_nb2%next\, \$1762_nb2%now\ : value(0 to 31) := (others => '0');
  signal \$1673_loop99401_arg%next\, \$1673_loop99401_arg%now\, 
         \$1831_loop99399_arg%next\, \$1831_loop99399_arg%now\, 
         \$1739_loop99401_arg%next\, \$1739_loop99401_arg%now\, 
         \$1607_loop99401_arg%next\, \$1607_loop99401_arg%now\, 
         \$1778_loop99400_arg%next\, \$1778_loop99400_arg%now\, 
         \$1619_loop99398_arg%next\, \$1619_loop99398_arg%now\, 
         \$1817_loop99398_arg%next\, \$1817_loop99398_arg%now\, 
         \$1805_loop99401_arg%next\, \$1805_loop99401_arg%now\, 
         \$1712_loop99400_arg%next\, \$1712_loop99400_arg%now\, 
         \$1699_loop99399_arg%next\, \$1699_loop99399_arg%now\, 
         \$1751_loop99398_arg%next\, \$1751_loop99398_arg%now\, 
         \$1765_loop99399_arg%next\, \$1765_loop99399_arg%now\, 
         \$1844_loop99400_arg%next\, \$1844_loop99400_arg%now\, 
         \$1633_loop99399_arg%next\, \$1633_loop99399_arg%now\, 
         \$1646_loop99400_arg%next\, \$1646_loop99400_arg%now\, 
         \$1685_loop99398_arg%next\, \$1685_loop99398_arg%now\ : value(0 to 415) := (others => '0');
  
  begin
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$$1209_src_write_request\ = '1' then
                    \$1209_src\(\$$1209_src_ptr_write\) <= \$$1209_src_write\;
                 end if;
                 \$$1209_src_value\ <= \$1209_src\(\$$1209_src_ptr\);
            end if;
        end process;
    
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$$1216_dst_write_request\ = '1' then
                    \$1216_dst\(\$$1216_dst_ptr_write\) <= \$$1216_dst_write\;
                 end if;
                 \$$1216_dst_value\ <= \$1216_dst\(\$$1216_dst_ptr\);
            end if;
        end process;
    
    process (clk)
            begin
            if rising_edge(clk) then
                 if \$$1217_r_write_request\ = '1' then
                    \$1217_r\(\$$1217_r_ptr_write\) <= \$$1217_r_write\;
                 end if;
                 \$$1217_r_value\ <= \$1217_r\(\$$1217_r_ptr\);
            end if;
        end process;
    
    process (reset,clk)
      begin
      if reset = '1' then
        \rdy569%now\ <= (others => '0');
        \$1737%now\ <= (others => '0');
        \$1646_loop99400_id%now\ <= (others => '0');
        \$1685_loop99398_arg%now\ <= (others => '0');
        \$v511%now\ <= (others => '0');
        \$1664%now\ <= (others => '0');
        \$1744%now\ <= (others => '0');
        \$1682%now\ <= (others => '0');
        \$1762_nb2%now\ <= (others => '0');
        \$v596%now\ <= (others => '0');
        \$1577_o%now\ <= (others => '0');
        \$v447%now\ <= (others => '0');
        \$1666%now\ <= (others => '0');
        \$1834%now\ <= (others => '0');
        \$1683%now\ <= (others => '0');
        \$1633_loop99399_result%now\ <= (others => '0');
        \$1637%now\ <= (others => '0');
        \$1646_loop99400_arg%now\ <= (others => '0');
        \$1803%now\ <= (others => '0');
        \$1797_n%now\ <= (others => '0');
        \$1698%now\ <= (others => '0');
        \$1735%now\ <= (others => '0');
        \$1730%now\ <= (others => '0');
        \$1685_loop99398_result%now\ <= (others => '0');
        \$v561%now\ <= (others => '0');
        \$1756%now\ <= (others => '0');
        \$1765_loop99399_id%now\ <= (others => '0');
        \$v579%now\ <= (others => '0');
        \$v557%now\ <= (others => '0');
        \$1719%now\ <= (others => '0');
        \$v413%now\ <= (others => '0');
        \$1811%now\ <= (others => '0');
        \$1703%now\ <= (others => '0');
        \$1821%now\ <= (others => '0');
        \$1640%now\ <= (others => '0');
        \$1633_loop99399_arg%now\ <= (others => '0');
        \$v553%now\ <= (others => '0');
        \$1645%now\ <= (others => '0');
        \$1627%now\ <= (others => '0');
        \$1613%now\ <= (others => '0');
        \$1712_loop99400_id%now\ <= (others => '0');
        \$1578%now\ <= (others => '0');
        \$1707%now\ <= (others => '0');
        \$1814%now\ <= (others => '0');
        \result574%now\ <= (others => '0');
        \$1755%now\ <= (others => '0');
        \$1677%now\ <= (others => '0');
        \result460%now\ <= (others => '0');
        \$1638%now\ <= (others => '0');
        \$v512%now\ <= (others => '0');
        \result502%now\ <= (others => '0');
        \$1815%now\ <= (others => '0');
        \$1771%now\ <= (others => '0');
        \$1684_nb2%now\ <= (others => '0');
        \$1660_id%now\ <= (others => '0');
        \$v550%now\ <= (others => '0');
        \result544%now\ <= (others => '0');
        \$v507%now\ <= (others => '0');
        \$v406%now\ <= (others => '0');
        \$1844_loop99400_arg%now\ <= (others => '0');
        \$1816_nb2%now\ <= (others => '0');
        \$1791_i%now\ <= (others => '0');
        \$1843%now\ <= (others => '0');
        \$1817_loop99398_id%now\ <= (others => '0');
        \result484%now\ <= (others => '0');
        \$1628%now\ <= (others => '0');
        \result403%now\ <= (others => '0');
        \$v513%now\ <= (others => '0');
        \$1639%now\ <= (others => '0');
        \$v540%now\ <= (others => '0');
        \$v517%now\ <= (others => '0');
        \$1665_n%now\ <= (others => '0');
        \$v543%now\ <= (others => '0');
        \rdy491%now\ <= (others => '0');
        \rdy408%now\ <= (others => '0');
        \$1597_i%now\ <= (others => '0');
        \$1860%now\ <= (others => '0');
        \$1852%now\ <= (others => '0');
        \$1787%now\ <= (others => '0');
        \$1705%now\ <= (others => '0');
        \$1593_i%now\ <= (others => '0');
        \$1853%now\ <= (others => '0');
        \$1831_loop99399_result%now\ <= (others => '0');
        \$1765_loop99399_arg%now\ <= (others => '0');
        \$1710_nb2%now\ <= (others => '0');
        \$v581%now\ <= (others => '0');
        \$v427%now\ <= (others => '0');
        \$1732%now\ <= (others => '0');
        \$1585%now\ <= (others => '0');
        \$1736%now\ <= (others => '0');
        \$1594_id%now\ <= (others => '0');
        \$v471%now\ <= (others => '0');
        \$1678%now\ <= (others => '0');
        \$1592%now\ <= (others => '0');
        \$1726_id%now\ <= (others => '0');
        \$1697%now\ <= (others => '0');
        \$1594_result%now\ <= (others => '0');
        \$1850%now\ <= (others => '0');
        \$v425%now\ <= (others => '0');
        \$1603%now\ <= (others => '0');
        \$1681%now\ <= (others => '0');
        \$1725_i%now\ <= (others => '0');
        \result568%now\ <= (others => '0');
        \$1672%now\ <= (others => '0');
        \$1790%now\ <= (others => '0');
        \$1782%now\ <= (others => '0');
        \$1649%now\ <= (others => '0');
        \$1623%now\ <= (others => '0');
        \$1856%now\ <= (others => '0');
        \$1825%now\ <= (others => '0');
        \$v539%now\ <= (others => '0');
        \$1622%now\ <= (others => '0');
        \$v497%now\ <= (others => '0');
        \$1583%now\ <= (others => '0');
        \$1792_id%now\ <= (others => '0');
        \$1751_loop99398_result%now\ <= (others => '0');
        \$1751_loop99398_arg%now\ <= (others => '0');
        \$1611%now\ <= (others => '0');
        \$1734%now\ <= (others => '0');
        \$1724%now\ <= (others => '0');
        \$v469%now\ <= (others => '0');
        \$v470%now\ <= (others => '0');
        \$1669%now\ <= (others => '0');
        \$1835%now\ <= (others => '0');
        \$1693%now\ <= (others => '0');
        \$v395%now\ <= (others => '0');
        \$v431%now\ <= (others => '0');
        \$v559%now\ <= (others => '0');
        \$v433%now\ <= (others => '0');
        \$v495%now\ <= (others => '0');
        \$1673_loop99401_id%now\ <= (others => '0');
        \$1691%now\ <= (others => '0');
        \$v481%now\ <= (others => '0');
        \$1716%now\ <= (others => '0');
        \$1601%now\ <= (others => '0');
        \$1702%now\ <= (others => '0');
        \$v432%now\ <= (others => '0');
        \$1625%now\ <= (others => '0');
        \$1857_id%now\ <= (others => '0');
        \$1745%now\ <= (others => '0');
        \$1685_loop99398_id%now\ <= (others => '0');
        \$1848%now\ <= (others => '0');
        \$1830%now\ <= (others => '0');
        \$1742%now\ <= (others => '0');
        \result418%now\ <= (others => '0');
        \$1692%now\ <= (others => '0');
        \$1581%now\ <= (others => '0');
        \$1591_x%now\ <= (others => '0');
        \$1776_nb2%now\ <= (others => '0');
        \$1676%now\ <= (others => '0');
        \$v590%now\ <= (others => '0');
        \$v478%now\ <= (others => '0');
        \$1670%now\ <= (others => '0');
        \$1739_loop99401_id%now\ <= (others => '0');
        \$1653%now\ <= (others => '0');
        \$1699_loop99399_arg%now\ <= (others => '0');
        \$1587%now\ <= (others => '0');
        \$v516%now\ <= (others => '0');
        \$1837%now\ <= (others => '0');
        \$v428%now\ <= (others => '0');
        \$v473%now\ <= (others => '0');
        \$v467%now\ <= (others => '0');
        \$1712_loop99400_arg%now\ <= (others => '0');
        \$1607_loop99401_id%now\ <= (others => '0');
        \$1715%now\ <= (others => '0');
        \$v466%now\ <= (others => '0');
        \$v562%now\ <= (others => '0');
        \$v501%now\ <= (others => '0');
        \$v593%now\ <= (others => '0');
        \$1659_i%now\ <= (others => '0');
        \$1827%now\ <= (others => '0');
        \$1617%now\ <= (others => '0');
        \$1750_nb2%now\ <= (others => '0');
        \$v435%now\ <= (others => '0');
        \$1851%now\ <= (others => '0');
        \$1743%now\ <= (others => '0');
        \$v573%now\ <= (others => '0');
        \$1788%now\ <= (others => '0');
        \rdy419%now\ <= (others => '0');
        \$v520%now\ <= (others => '0');
        \$1854%now\ <= (others => '0');
        \$v565%now\ <= (others => '0');
        \$1805_loop99401_arg%now\ <= (others => '0');
        \$1781%now\ <= (others => '0');
        \rdy461%now\ <= (others => '0');
        \rdy404%now\ <= (others => '0');
        \result448%now\ <= (others => '0');
        \$v429%now\ <= (others => '0');
        \$1694%now\ <= (others => '0');
        \$1840%now\ <= (others => '0');
        \$1775%now\ <= (others => '0');
        \$1629%now\ <= (others => '0');
        \$1712_loop99400_result%now\ <= (others => '0');
        \$v480%now\ <= (others => '0');
        \rdy527%now\ <= (others => '0');
        \$v509%now\ <= (others => '0');
        \rdy485%now\ <= (others => '0');
        \$1778_loop99400_id%now\ <= (others => '0');
        \$1588_id%now\ <= (others => '0');
        \$1841%now\ <= (others => '0');
        \$1817_loop99398_arg%now\ <= (others => '0');
        \$v459%now\ <= (others => '0');
        \$1792_result%now\ <= (others => '0');
        \$1768%now\ <= (others => '0');
        \$1632%now\ <= (others => '0');
        \$v521%now\ <= (others => '0');
        \$v476%now\ <= (others => '0');
        \$1598%now\ <= (others => '0');
        \$1657_nb2%now\ <= (others => '0');
        \$1644_nb2%now\ <= (others => '0');
        \$1696_nb2%now\ <= (others => '0');
        \$v438%now\ <= (others => '0');
        \$v555%now\ <= (others => '0');
        \$1718%now\ <= (others => '0');
        \$1796%now\ <= (others => '0');
        \$1844_loop99400_id%now\ <= (others => '0');
        \$v424%now\ <= (others => '0');
        \$1584%now\ <= (others => '0');
        \$1855_nb2%now\ <= (others => '0');
        \$v456%now\ <= (others => '0');
        \$1619_loop99398_id%now\ <= (others => '0');
        \$1817_loop99398_result%now\ <= (others => '0');
        \$1642%now\ <= (others => '0');
        \$1619_loop99398_arg%now\ <= (others => '0');
        \$v426%now\ <= (others => '0');
        \$v397%now\ <= (others => '0');
        \$1689%now\ <= (others => '0');
        \$1847%now\ <= (others => '0');
        \$1679%now\ <= (others => '0');
        \result442%now\ <= (others => '0');
        \$1844_loop99400_result%now\ <= (others => '0');
        \$v537%now\ <= (others => '0');
        \$1783%now\ <= (others => '0');
        \$v489%now\ <= (others => '0');
        \$1809%now\ <= (others => '0');
        \$1849%now\ <= (others => '0');
        \$1607_loop99401_result%now\ <= (others => '0');
        \$v436%now\ <= (others => '0');
        \$1826%now\ <= (others => '0');
        \$v472%now\ <= (others => '0');
        \$v434%now\ <= (others => '0');
        \$1602%now\ <= (others => '0');
        \$1792_arg%now\ <= (others => '0');
        \result407%now\ <= (others => '0');
        \$1778_loop99400_result%now\ <= (others => '0');
        \$1761%now\ <= (others => '0');
        \$1708%now\ <= (others => '0');
        \$1599_n%now\ <= (others => '0');
        \$v479%now\ <= (others => '0');
        \$1748%now\ <= (others => '0');
        \$1800%now\ <= (others => '0');
        \$1823%now\ <= (others => '0');
        \$v554%now\ <= (others => '0');
        \$1726_result%now\ <= (others => '0');
        \$1626%now\ <= (others => '0');
        \$v552%now\ <= (others => '0');
        \$1824%now\ <= (others => '0');
        \$1695%now\ <= (others => '0');
        \$1699_loop99399_id%now\ <= (others => '0');
        \$1739_loop99401_result%now\ <= (others => '0');
        \$1747%now\ <= (others => '0');
        \$v498%now\ <= (others => '0');
        \$1650%now\ <= (others => '0');
        \$1624%now\ <= (others => '0');
        \$1839%now\ <= (others => '0');
        \$1651%now\ <= (others => '0');
        \$1667%now\ <= (others => '0');
        \$1673_loop99401_result%now\ <= (others => '0');
        \$1652%now\ <= (others => '0');
        \$1646_loop99400_result%now\ <= (others => '0');
        \$1802%now\ <= (others => '0');
        \$1777%now\ <= (others => '0');
        \$1671%now\ <= (others => '0');
        \$1757%now\ <= (others => '0');
        \$v453%now\ <= (others => '0');
        \$1720%now\ <= (others => '0');
        \$v563%now\ <= (others => '0');
        \$1749%now\ <= (others => '0');
        \$v549%now\ <= (others => '0');
        \$v585%now\ <= (others => '0');
        \$v423%now\ <= (others => '0');
        \$1805_loop99401_id%now\ <= (others => '0');
        \$1699_loop99399_result%now\ <= (others => '0');
        \$1842_nb2%now\ <= (others => '0');
        \$1774%now\ <= (others => '0');
        \$1723_nb2%now\ <= (others => '0');
        \$1633_loop99399_id%now\ <= (others => '0');
        \$1612%now\ <= (others => '0');
        \$1829%now\ <= (others => '0');
        \$1785%now\ <= (others => '0');
        \$1733%now\ <= (others => '0');
        \$1773%now\ <= (others => '0');
        \$v515%now\ <= (others => '0');
        \$v439%now\ <= (others => '0');
        \$v551%now\ <= (others => '0');
        \$1688%now\ <= (others => '0');
        \$1582%now\ <= (others => '0');
        \$v430%now\ <= (others => '0');
        \rdy545%now\ <= (others => '0');
        \$1822%now\ <= (others => '0');
        \$1654%now\ <= (others => '0');
        \$1786%now\ <= (others => '0');
        \$1828_nb2%now\ <= (others => '0');
        \$1798%now\ <= (others => '0');
        \$1778_loop99400_arg%now\ <= (others => '0');
        \$1857_result%now\ <= (others => '0');
        \$1660_arg%now\ <= (others => '0');
        \$1641%now\ <= (others => '0');
        \$1769%now\ <= (others => '0');
        \rdy449%now\ <= (others => '0');
        \$1857_arg%now\ <= (others => '0');
        \$1726_arg%now\ <= (others => '0');
        \$1610%now\ <= (others => '0');
        \$1804%now\ <= (others => '0');
        \$1754%now\ <= (others => '0');
        \$1759%now\ <= (others => '0');
        \$v465%now\ <= (others => '0');
        \$v531%now\ <= (others => '0');
        \$v508%now\ <= (others => '0');
        \$1643%now\ <= (others => '0');
        \result490%now\ <= (others => '0');
        \$v564%now\ <= (others => '0');
        \$1656%now\ <= (others => '0');
        \$v437%now\ <= (others => '0');
        \$1586%now\ <= (others => '0');
        \$1760%now\ <= (others => '0');
        \$1813%now\ <= (others => '0');
        \$1721%now\ <= (others => '0');
        \$1680%now\ <= (others => '0');
        \$v522%now\ <= (others => '0');
        \$1668%now\ <= (others => '0');
        \$1831_loop99399_id%now\ <= (others => '0');
        \result526%now\ <= (others => '0');
        \$1746%now\ <= (others => '0');
        \$v560%now\ <= (others => '0');
        \rdy443%now\ <= (others => '0');
        \$v475%now\ <= (others => '0');
        \$1588_result%now\ <= (others => '0');
        \$v477%now\ <= (others => '0');
        \$1607_loop99401_arg%now\ <= (others => '0');
        \$1631%now\ <= (others => '0');
        \$v582%now\ <= (others => '0');
        \$v514%now\ <= (others => '0');
        \$1772%now\ <= (others => '0');
        \$1739_loop99401_arg%now\ <= (others => '0');
        \$v455%now\ <= (others => '0');
        \$1580_led%now\ <= (others => '0');
        \$v587%now\ <= (others => '0');
        \$1605%now\ <= (others => '0');
        \$1820%now\ <= (others => '0');
        \$v468%now\ <= (others => '0');
        \rdy575%now\ <= (others => '0');
        \$1801%now\ <= (others => '0');
        \$1660_result%now\ <= (others => '0');
        \$v556%now\ <= (others => '0');
        \$1861%now\ <= (others => '0');
        \$1764%now\ <= (others => '0');
        \$1836%now\ <= (others => '0');
        \$1838%now\ <= (others => '0');
        \$v558%now\ <= (others => '0');
        \$1738%now\ <= (others => '0');
        \$1630_nb2%now\ <= (others => '0');
        \$1579%now\ <= (others => '0');
        \$1805_loop99401_result%now\ <= (others => '0');
        \$1729_i%now\ <= (others => '0');
        \$1751_loop99398_id%now\ <= (others => '0');
        \$1722%now\ <= (others => '0');
        \$1618_nb2%now\ <= (others => '0');
        \$1795_i%now\ <= (others => '0');
        \$1758%now\ <= (others => '0');
        \$1658%now\ <= (others => '0');
        \$v519%now\ <= (others => '0');
        \$1784%now\ <= (others => '0');
        \$1763%now\ <= (others => '0');
        \$1588_arg%now\ <= (others => '0');
        \$1616%now\ <= (others => '0');
        \$1808%now\ <= (others => '0');
        \result532%now\ <= (others => '0');
        \$1655%now\ <= (others => '0');
        \$v594%now\ <= (others => '0');
        \rdy533%now\ <= (others => '0');
        \$1765_loop99399_result%now\ <= (others => '0');
        \$v523%now\ <= (others => '0');
        \$1604%now\ <= (others => '0');
        \$1711%now\ <= (others => '0');
        \$1663_i%now\ <= (others => '0');
        \$1636%now\ <= (others => '0');
        \$1799%now\ <= (others => '0');
        \$1810%now\ <= (others => '0');
        \$1831_loop99399_arg%now\ <= (others => '0');
        \$1731_n%now\ <= (others => '0');
        \$v474%now\ <= (others => '0');
        \$v510%now\ <= (others => '0');
        \$1594_arg%now\ <= (others => '0');
        \$1615%now\ <= (others => '0');
        \$v518%now\ <= (others => '0');
        \$1717%now\ <= (others => '0');
        \$1706%now\ <= (others => '0');
        \$1606%now\ <= (others => '0');
        \$1789_nb2%now\ <= (others => '0');
        \$1600%now\ <= (others => '0');
        \$1770%now\ <= (others => '0');
        \$1709%now\ <= (others => '0');
        \$1673_loop99401_arg%now\ <= (others => '0');
        \$1704%now\ <= (others => '0');
        \$1690%now\ <= (others => '0');
        \$1619_loop99398_result%now\ <= (others => '0');
        \rdy503%now\ <= (others => '0');
        \$1812%now\ <= (others => '0');
        \$1614%now\ <= (others => '0');
        \$v412%now\ <= (others => '0');
        \$$1209_src_lock%now\ <= (others => '0');
        \$$1216_dst_lock%now\ <= (others => '0');
        \$$1217_r_lock%now\ <= (others => '0');
        \state%now\ <= idle405;
        \state_var609%now\ <= idle444;
        \state_var608%now\ <= idle450;
        \state_var607%now\ <= idle420;
        \state_var606%now\ <= idle486;
        \state_var605%now\ <= idle492;
        \state_var604%now\ <= idle462;
        \state_var603%now\ <= idle528;
        \state_var602%now\ <= idle534;
        \state_var601%now\ <= idle504;
        \state_var600%now\ <= idle570;
        \state_var599%now\ <= idle576;
        \state_var598%now\ <= idle546;
        \state_var597%now\ <= idle409;
      elsif (rising_edge(clk)) then
        \rdy569%now\ <= \rdy569%next\;
        \$1737%now\ <= \$1737%next\;
        \$1646_loop99400_id%now\ <= \$1646_loop99400_id%next\;
        \$1685_loop99398_arg%now\ <= \$1685_loop99398_arg%next\;
        \$v511%now\ <= \$v511%next\;
        \$1664%now\ <= \$1664%next\;
        \$1744%now\ <= \$1744%next\;
        \$1682%now\ <= \$1682%next\;
        \$1762_nb2%now\ <= \$1762_nb2%next\;
        \$v596%now\ <= \$v596%next\;
        \$1577_o%now\ <= \$1577_o%next\;
        \$v447%now\ <= \$v447%next\;
        \$1666%now\ <= \$1666%next\;
        \$1834%now\ <= \$1834%next\;
        \$1683%now\ <= \$1683%next\;
        \$1633_loop99399_result%now\ <= \$1633_loop99399_result%next\;
        \$1637%now\ <= \$1637%next\;
        \$1646_loop99400_arg%now\ <= \$1646_loop99400_arg%next\;
        \$1803%now\ <= \$1803%next\;
        \$1797_n%now\ <= \$1797_n%next\;
        \$1698%now\ <= \$1698%next\;
        \$1735%now\ <= \$1735%next\;
        \$1730%now\ <= \$1730%next\;
        \$1685_loop99398_result%now\ <= \$1685_loop99398_result%next\;
        \$v561%now\ <= \$v561%next\;
        \$1756%now\ <= \$1756%next\;
        \$1765_loop99399_id%now\ <= \$1765_loop99399_id%next\;
        \$v579%now\ <= \$v579%next\;
        \$v557%now\ <= \$v557%next\;
        \$1719%now\ <= \$1719%next\;
        \$v413%now\ <= \$v413%next\;
        \$1811%now\ <= \$1811%next\;
        \$1703%now\ <= \$1703%next\;
        \$1821%now\ <= \$1821%next\;
        \$1640%now\ <= \$1640%next\;
        \$1633_loop99399_arg%now\ <= \$1633_loop99399_arg%next\;
        \$v553%now\ <= \$v553%next\;
        \$1645%now\ <= \$1645%next\;
        \$1627%now\ <= \$1627%next\;
        \$1613%now\ <= \$1613%next\;
        \$1712_loop99400_id%now\ <= \$1712_loop99400_id%next\;
        \$1578%now\ <= \$1578%next\;
        \$1707%now\ <= \$1707%next\;
        \$1814%now\ <= \$1814%next\;
        \result574%now\ <= \result574%next\;
        \$1755%now\ <= \$1755%next\;
        \$1677%now\ <= \$1677%next\;
        \result460%now\ <= \result460%next\;
        \$1638%now\ <= \$1638%next\;
        \$v512%now\ <= \$v512%next\;
        \result502%now\ <= \result502%next\;
        \$1815%now\ <= \$1815%next\;
        \$1771%now\ <= \$1771%next\;
        \$1684_nb2%now\ <= \$1684_nb2%next\;
        \$1660_id%now\ <= \$1660_id%next\;
        \$v550%now\ <= \$v550%next\;
        \result544%now\ <= \result544%next\;
        \$v507%now\ <= \$v507%next\;
        \$v406%now\ <= \$v406%next\;
        \$1844_loop99400_arg%now\ <= \$1844_loop99400_arg%next\;
        \$1816_nb2%now\ <= \$1816_nb2%next\;
        \$1791_i%now\ <= \$1791_i%next\;
        \$1843%now\ <= \$1843%next\;
        \$1817_loop99398_id%now\ <= \$1817_loop99398_id%next\;
        \result484%now\ <= \result484%next\;
        \$1628%now\ <= \$1628%next\;
        \result403%now\ <= \result403%next\;
        \$v513%now\ <= \$v513%next\;
        \$1639%now\ <= \$1639%next\;
        \$v540%now\ <= \$v540%next\;
        \$v517%now\ <= \$v517%next\;
        \$1665_n%now\ <= \$1665_n%next\;
        \$v543%now\ <= \$v543%next\;
        \rdy491%now\ <= \rdy491%next\;
        \rdy408%now\ <= \rdy408%next\;
        \$1597_i%now\ <= \$1597_i%next\;
        \$1860%now\ <= \$1860%next\;
        \$1852%now\ <= \$1852%next\;
        \$1787%now\ <= \$1787%next\;
        \$1705%now\ <= \$1705%next\;
        \$1593_i%now\ <= \$1593_i%next\;
        \$1853%now\ <= \$1853%next\;
        \$1831_loop99399_result%now\ <= \$1831_loop99399_result%next\;
        \$1765_loop99399_arg%now\ <= \$1765_loop99399_arg%next\;
        \$1710_nb2%now\ <= \$1710_nb2%next\;
        \$v581%now\ <= \$v581%next\;
        \$v427%now\ <= \$v427%next\;
        \$1732%now\ <= \$1732%next\;
        \$1585%now\ <= \$1585%next\;
        \$1736%now\ <= \$1736%next\;
        \$1594_id%now\ <= \$1594_id%next\;
        \$v471%now\ <= \$v471%next\;
        \$1678%now\ <= \$1678%next\;
        \$1592%now\ <= \$1592%next\;
        \$1726_id%now\ <= \$1726_id%next\;
        \$1697%now\ <= \$1697%next\;
        \$1594_result%now\ <= \$1594_result%next\;
        \$1850%now\ <= \$1850%next\;
        \$v425%now\ <= \$v425%next\;
        \$1603%now\ <= \$1603%next\;
        \$1681%now\ <= \$1681%next\;
        \$1725_i%now\ <= \$1725_i%next\;
        \result568%now\ <= \result568%next\;
        \$1672%now\ <= \$1672%next\;
        \$1790%now\ <= \$1790%next\;
        \$1782%now\ <= \$1782%next\;
        \$1649%now\ <= \$1649%next\;
        \$1623%now\ <= \$1623%next\;
        \$1856%now\ <= \$1856%next\;
        \$1825%now\ <= \$1825%next\;
        \$v539%now\ <= \$v539%next\;
        \$1622%now\ <= \$1622%next\;
        \$v497%now\ <= \$v497%next\;
        \$1583%now\ <= \$1583%next\;
        \$1792_id%now\ <= \$1792_id%next\;
        \$1751_loop99398_result%now\ <= \$1751_loop99398_result%next\;
        \$1751_loop99398_arg%now\ <= \$1751_loop99398_arg%next\;
        \$1611%now\ <= \$1611%next\;
        \$1734%now\ <= \$1734%next\;
        \$1724%now\ <= \$1724%next\;
        \$v469%now\ <= \$v469%next\;
        \$v470%now\ <= \$v470%next\;
        \$1669%now\ <= \$1669%next\;
        \$1835%now\ <= \$1835%next\;
        \$1693%now\ <= \$1693%next\;
        \$v395%now\ <= \$v395%next\;
        \$v431%now\ <= \$v431%next\;
        \$v559%now\ <= \$v559%next\;
        \$v433%now\ <= \$v433%next\;
        \$v495%now\ <= \$v495%next\;
        \$1673_loop99401_id%now\ <= \$1673_loop99401_id%next\;
        \$1691%now\ <= \$1691%next\;
        \$v481%now\ <= \$v481%next\;
        \$1716%now\ <= \$1716%next\;
        \$1601%now\ <= \$1601%next\;
        \$1702%now\ <= \$1702%next\;
        \$v432%now\ <= \$v432%next\;
        \$1625%now\ <= \$1625%next\;
        \$1857_id%now\ <= \$1857_id%next\;
        \$1745%now\ <= \$1745%next\;
        \$1685_loop99398_id%now\ <= \$1685_loop99398_id%next\;
        \$1848%now\ <= \$1848%next\;
        \$1830%now\ <= \$1830%next\;
        \$1742%now\ <= \$1742%next\;
        \result418%now\ <= \result418%next\;
        \$1692%now\ <= \$1692%next\;
        \$1581%now\ <= \$1581%next\;
        \$1591_x%now\ <= \$1591_x%next\;
        \$1776_nb2%now\ <= \$1776_nb2%next\;
        \$1676%now\ <= \$1676%next\;
        \$v590%now\ <= \$v590%next\;
        \$v478%now\ <= \$v478%next\;
        \$1670%now\ <= \$1670%next\;
        \$1739_loop99401_id%now\ <= \$1739_loop99401_id%next\;
        \$1653%now\ <= \$1653%next\;
        \$1699_loop99399_arg%now\ <= \$1699_loop99399_arg%next\;
        \$1587%now\ <= \$1587%next\;
        \$v516%now\ <= \$v516%next\;
        \$1837%now\ <= \$1837%next\;
        \$v428%now\ <= \$v428%next\;
        \$v473%now\ <= \$v473%next\;
        \$v467%now\ <= \$v467%next\;
        \$1712_loop99400_arg%now\ <= \$1712_loop99400_arg%next\;
        \$1607_loop99401_id%now\ <= \$1607_loop99401_id%next\;
        \$1715%now\ <= \$1715%next\;
        \$v466%now\ <= \$v466%next\;
        \$v562%now\ <= \$v562%next\;
        \$v501%now\ <= \$v501%next\;
        \$v593%now\ <= \$v593%next\;
        \$1659_i%now\ <= \$1659_i%next\;
        \$1827%now\ <= \$1827%next\;
        \$1617%now\ <= \$1617%next\;
        \$1750_nb2%now\ <= \$1750_nb2%next\;
        \$v435%now\ <= \$v435%next\;
        \$1851%now\ <= \$1851%next\;
        \$1743%now\ <= \$1743%next\;
        \$v573%now\ <= \$v573%next\;
        \$1788%now\ <= \$1788%next\;
        \rdy419%now\ <= \rdy419%next\;
        \$v520%now\ <= \$v520%next\;
        \$1854%now\ <= \$1854%next\;
        \$v565%now\ <= \$v565%next\;
        \$1805_loop99401_arg%now\ <= \$1805_loop99401_arg%next\;
        \$1781%now\ <= \$1781%next\;
        \rdy461%now\ <= \rdy461%next\;
        \rdy404%now\ <= \rdy404%next\;
        \result448%now\ <= \result448%next\;
        \$v429%now\ <= \$v429%next\;
        \$1694%now\ <= \$1694%next\;
        \$1840%now\ <= \$1840%next\;
        \$1775%now\ <= \$1775%next\;
        \$1629%now\ <= \$1629%next\;
        \$1712_loop99400_result%now\ <= \$1712_loop99400_result%next\;
        \$v480%now\ <= \$v480%next\;
        \rdy527%now\ <= \rdy527%next\;
        \$v509%now\ <= \$v509%next\;
        \rdy485%now\ <= \rdy485%next\;
        \$1778_loop99400_id%now\ <= \$1778_loop99400_id%next\;
        \$1588_id%now\ <= \$1588_id%next\;
        \$1841%now\ <= \$1841%next\;
        \$1817_loop99398_arg%now\ <= \$1817_loop99398_arg%next\;
        \$v459%now\ <= \$v459%next\;
        \$1792_result%now\ <= \$1792_result%next\;
        \$1768%now\ <= \$1768%next\;
        \$1632%now\ <= \$1632%next\;
        \$v521%now\ <= \$v521%next\;
        \$v476%now\ <= \$v476%next\;
        \$1598%now\ <= \$1598%next\;
        \$1657_nb2%now\ <= \$1657_nb2%next\;
        \$1644_nb2%now\ <= \$1644_nb2%next\;
        \$1696_nb2%now\ <= \$1696_nb2%next\;
        \$v438%now\ <= \$v438%next\;
        \$v555%now\ <= \$v555%next\;
        \$1718%now\ <= \$1718%next\;
        \$1796%now\ <= \$1796%next\;
        \$1844_loop99400_id%now\ <= \$1844_loop99400_id%next\;
        \$v424%now\ <= \$v424%next\;
        \$1584%now\ <= \$1584%next\;
        \$1855_nb2%now\ <= \$1855_nb2%next\;
        \$v456%now\ <= \$v456%next\;
        \$1619_loop99398_id%now\ <= \$1619_loop99398_id%next\;
        \$1817_loop99398_result%now\ <= \$1817_loop99398_result%next\;
        \$1642%now\ <= \$1642%next\;
        \$1619_loop99398_arg%now\ <= \$1619_loop99398_arg%next\;
        \$v426%now\ <= \$v426%next\;
        \$v397%now\ <= \$v397%next\;
        \$1689%now\ <= \$1689%next\;
        \$1847%now\ <= \$1847%next\;
        \$1679%now\ <= \$1679%next\;
        \result442%now\ <= \result442%next\;
        \$1844_loop99400_result%now\ <= \$1844_loop99400_result%next\;
        \$v537%now\ <= \$v537%next\;
        \$1783%now\ <= \$1783%next\;
        \$v489%now\ <= \$v489%next\;
        \$1809%now\ <= \$1809%next\;
        \$1849%now\ <= \$1849%next\;
        \$1607_loop99401_result%now\ <= \$1607_loop99401_result%next\;
        \$v436%now\ <= \$v436%next\;
        \$1826%now\ <= \$1826%next\;
        \$v472%now\ <= \$v472%next\;
        \$v434%now\ <= \$v434%next\;
        \$1602%now\ <= \$1602%next\;
        \$1792_arg%now\ <= \$1792_arg%next\;
        \result407%now\ <= \result407%next\;
        \$1778_loop99400_result%now\ <= \$1778_loop99400_result%next\;
        \$1761%now\ <= \$1761%next\;
        \$1708%now\ <= \$1708%next\;
        \$1599_n%now\ <= \$1599_n%next\;
        \$v479%now\ <= \$v479%next\;
        \$1748%now\ <= \$1748%next\;
        \$1800%now\ <= \$1800%next\;
        \$1823%now\ <= \$1823%next\;
        \$v554%now\ <= \$v554%next\;
        \$1726_result%now\ <= \$1726_result%next\;
        \$1626%now\ <= \$1626%next\;
        \$v552%now\ <= \$v552%next\;
        \$1824%now\ <= \$1824%next\;
        \$1695%now\ <= \$1695%next\;
        \$1699_loop99399_id%now\ <= \$1699_loop99399_id%next\;
        \$1739_loop99401_result%now\ <= \$1739_loop99401_result%next\;
        \$1747%now\ <= \$1747%next\;
        \$v498%now\ <= \$v498%next\;
        \$1650%now\ <= \$1650%next\;
        \$1624%now\ <= \$1624%next\;
        \$1839%now\ <= \$1839%next\;
        \$1651%now\ <= \$1651%next\;
        \$1667%now\ <= \$1667%next\;
        \$1673_loop99401_result%now\ <= \$1673_loop99401_result%next\;
        \$1652%now\ <= \$1652%next\;
        \$1646_loop99400_result%now\ <= \$1646_loop99400_result%next\;
        \$1802%now\ <= \$1802%next\;
        \$1777%now\ <= \$1777%next\;
        \$1671%now\ <= \$1671%next\;
        \$1757%now\ <= \$1757%next\;
        \$v453%now\ <= \$v453%next\;
        \$1720%now\ <= \$1720%next\;
        \$v563%now\ <= \$v563%next\;
        \$1749%now\ <= \$1749%next\;
        \$v549%now\ <= \$v549%next\;
        \$v585%now\ <= \$v585%next\;
        \$v423%now\ <= \$v423%next\;
        \$1805_loop99401_id%now\ <= \$1805_loop99401_id%next\;
        \$1699_loop99399_result%now\ <= \$1699_loop99399_result%next\;
        \$1842_nb2%now\ <= \$1842_nb2%next\;
        \$1774%now\ <= \$1774%next\;
        \$1723_nb2%now\ <= \$1723_nb2%next\;
        \$1633_loop99399_id%now\ <= \$1633_loop99399_id%next\;
        \$1612%now\ <= \$1612%next\;
        \$1829%now\ <= \$1829%next\;
        \$1785%now\ <= \$1785%next\;
        \$1733%now\ <= \$1733%next\;
        \$1773%now\ <= \$1773%next\;
        \$v515%now\ <= \$v515%next\;
        \$v439%now\ <= \$v439%next\;
        \$v551%now\ <= \$v551%next\;
        \$1688%now\ <= \$1688%next\;
        \$1582%now\ <= \$1582%next\;
        \$v430%now\ <= \$v430%next\;
        \rdy545%now\ <= \rdy545%next\;
        \$1822%now\ <= \$1822%next\;
        \$1654%now\ <= \$1654%next\;
        \$1786%now\ <= \$1786%next\;
        \$1828_nb2%now\ <= \$1828_nb2%next\;
        \$1798%now\ <= \$1798%next\;
        \$1778_loop99400_arg%now\ <= \$1778_loop99400_arg%next\;
        \$1857_result%now\ <= \$1857_result%next\;
        \$1660_arg%now\ <= \$1660_arg%next\;
        \$1641%now\ <= \$1641%next\;
        \$1769%now\ <= \$1769%next\;
        \rdy449%now\ <= \rdy449%next\;
        \$1857_arg%now\ <= \$1857_arg%next\;
        \$1726_arg%now\ <= \$1726_arg%next\;
        \$1610%now\ <= \$1610%next\;
        \$1804%now\ <= \$1804%next\;
        \$1754%now\ <= \$1754%next\;
        \$1759%now\ <= \$1759%next\;
        \$v465%now\ <= \$v465%next\;
        \$v531%now\ <= \$v531%next\;
        \$v508%now\ <= \$v508%next\;
        \$1643%now\ <= \$1643%next\;
        \result490%now\ <= \result490%next\;
        \$v564%now\ <= \$v564%next\;
        \$1656%now\ <= \$1656%next\;
        \$v437%now\ <= \$v437%next\;
        \$1586%now\ <= \$1586%next\;
        \$1760%now\ <= \$1760%next\;
        \$1813%now\ <= \$1813%next\;
        \$1721%now\ <= \$1721%next\;
        \$1680%now\ <= \$1680%next\;
        \$v522%now\ <= \$v522%next\;
        \$1668%now\ <= \$1668%next\;
        \$1831_loop99399_id%now\ <= \$1831_loop99399_id%next\;
        \result526%now\ <= \result526%next\;
        \$1746%now\ <= \$1746%next\;
        \$v560%now\ <= \$v560%next\;
        \rdy443%now\ <= \rdy443%next\;
        \$v475%now\ <= \$v475%next\;
        \$1588_result%now\ <= \$1588_result%next\;
        \$v477%now\ <= \$v477%next\;
        \$1607_loop99401_arg%now\ <= \$1607_loop99401_arg%next\;
        \$1631%now\ <= \$1631%next\;
        \$v582%now\ <= \$v582%next\;
        \$v514%now\ <= \$v514%next\;
        \$1772%now\ <= \$1772%next\;
        \$1739_loop99401_arg%now\ <= \$1739_loop99401_arg%next\;
        \$v455%now\ <= \$v455%next\;
        \$1580_led%now\ <= \$1580_led%next\;
        \$v587%now\ <= \$v587%next\;
        \$1605%now\ <= \$1605%next\;
        \$1820%now\ <= \$1820%next\;
        \$v468%now\ <= \$v468%next\;
        \rdy575%now\ <= \rdy575%next\;
        \$1801%now\ <= \$1801%next\;
        \$1660_result%now\ <= \$1660_result%next\;
        \$v556%now\ <= \$v556%next\;
        \$1861%now\ <= \$1861%next\;
        \$1764%now\ <= \$1764%next\;
        \$1836%now\ <= \$1836%next\;
        \$1838%now\ <= \$1838%next\;
        \$v558%now\ <= \$v558%next\;
        \$1738%now\ <= \$1738%next\;
        \$1630_nb2%now\ <= \$1630_nb2%next\;
        \$1579%now\ <= \$1579%next\;
        \$1805_loop99401_result%now\ <= \$1805_loop99401_result%next\;
        \$1729_i%now\ <= \$1729_i%next\;
        \$1751_loop99398_id%now\ <= \$1751_loop99398_id%next\;
        \$1722%now\ <= \$1722%next\;
        \$1618_nb2%now\ <= \$1618_nb2%next\;
        \$1795_i%now\ <= \$1795_i%next\;
        \$1758%now\ <= \$1758%next\;
        \$1658%now\ <= \$1658%next\;
        \$v519%now\ <= \$v519%next\;
        \$1784%now\ <= \$1784%next\;
        \$1763%now\ <= \$1763%next\;
        \$1588_arg%now\ <= \$1588_arg%next\;
        \$1616%now\ <= \$1616%next\;
        \$1808%now\ <= \$1808%next\;
        \result532%now\ <= \result532%next\;
        \$1655%now\ <= \$1655%next\;
        \$v594%now\ <= \$v594%next\;
        \rdy533%now\ <= \rdy533%next\;
        \$1765_loop99399_result%now\ <= \$1765_loop99399_result%next\;
        \$v523%now\ <= \$v523%next\;
        \$1604%now\ <= \$1604%next\;
        \$1711%now\ <= \$1711%next\;
        \$1663_i%now\ <= \$1663_i%next\;
        \$1636%now\ <= \$1636%next\;
        \$1799%now\ <= \$1799%next\;
        \$1810%now\ <= \$1810%next\;
        \$1831_loop99399_arg%now\ <= \$1831_loop99399_arg%next\;
        \$1731_n%now\ <= \$1731_n%next\;
        \$v474%now\ <= \$v474%next\;
        \$v510%now\ <= \$v510%next\;
        \$1594_arg%now\ <= \$1594_arg%next\;
        \$1615%now\ <= \$1615%next\;
        \$v518%now\ <= \$v518%next\;
        \$1717%now\ <= \$1717%next\;
        \$1706%now\ <= \$1706%next\;
        \$1606%now\ <= \$1606%next\;
        \$1789_nb2%now\ <= \$1789_nb2%next\;
        \$1600%now\ <= \$1600%next\;
        \$1770%now\ <= \$1770%next\;
        \$1709%now\ <= \$1709%next\;
        \$1673_loop99401_arg%now\ <= \$1673_loop99401_arg%next\;
        \$1704%now\ <= \$1704%next\;
        \$1690%now\ <= \$1690%next\;
        \$1619_loop99398_result%now\ <= \$1619_loop99398_result%next\;
        \rdy503%now\ <= \rdy503%next\;
        \$1812%now\ <= \$1812%next\;
        \$1614%now\ <= \$1614%next\;
        \$v412%now\ <= \$v412%next\;
        \$$1209_src_lock%now\ <= \$$1209_src_lock%next\;
        \$$1216_dst_lock%now\ <= \$$1216_dst_lock%next\;
        \$$1217_r_lock%now\ <= \$$1217_r_lock%next\;
        \state_var609%now\ <= \state_var609%next\;
        \state_var608%now\ <= \state_var608%next\;
        \state_var607%now\ <= \state_var607%next\;
        \state_var606%now\ <= \state_var606%next\;
        \state_var605%now\ <= \state_var605%next\;
        \state_var604%now\ <= \state_var604%next\;
        \state_var603%now\ <= \state_var603%next\;
        \state_var602%now\ <= \state_var602%next\;
        \state_var601%now\ <= \state_var601%next\;
        \state_var600%now\ <= \state_var600%next\;
        \state_var599%now\ <= \state_var599%next\;
        \state_var598%now\ <= \state_var598%next\;
        \state_var597%now\ <= \state_var597%next\;
        \state%now\ <= \state%next\;
      end if;
    end process;
      
      process(argument,\state%now\, clk,\state_var609%now\,\state_var608%now\,\state_var607%now\,\state_var606%now\,\state_var605%now\,\state_var604%now\,\state_var603%now\,\state_var602%now\,\state_var601%now\,\state_var600%now\,\state_var599%now\,\state_var598%now\,\state_var597%now\, \$$1209_src_value\, \$$1216_dst_value\, \$$1217_r_value\, \rdy569%now\, \$1737%now\, \$1646_loop99400_id%now\, \$1685_loop99398_arg%now\, \$v511%now\, \$1664%now\, \$1744%now\, \$1682%now\, \$1762_nb2%now\, \$v596%now\, \$1577_o%now\, \$v447%now\, \$1666%now\, \$1834%now\, \$1683%now\, \$1633_loop99399_result%now\, \$1637%now\, \$1646_loop99400_arg%now\, \$1803%now\, \$1797_n%now\, \$1698%now\, \$1735%now\, \$1730%now\, \$1685_loop99398_result%now\, \$v561%now\, \$1756%now\, \$1765_loop99399_id%now\, \$v579%now\, \$v557%now\, \$1719%now\, \$v413%now\, \$1811%now\, \$1703%now\, \$1821%now\, \$1640%now\, \$1633_loop99399_arg%now\, \$v553%now\, \$1645%now\, \$1627%now\, \$1613%now\, \$1712_loop99400_id%now\, \$1578%now\, \$1707%now\, \$1814%now\, \result574%now\, \$1755%now\, \$1677%now\, \result460%now\, \$1638%now\, \$v512%now\, \result502%now\, \$1815%now\, \$1771%now\, \$1684_nb2%now\, \$1660_id%now\, \$v550%now\, \result544%now\, \$v507%now\, \$v406%now\, \$1844_loop99400_arg%now\, \$1816_nb2%now\, \$1791_i%now\, \$1843%now\, \$1817_loop99398_id%now\, \result484%now\, \$1628%now\, \result403%now\, \$v513%now\, \$1639%now\, \$v540%now\, \$v517%now\, \$1665_n%now\, \$v543%now\, \rdy491%now\, \rdy408%now\, \$1597_i%now\, \$1860%now\, \$1852%now\, \$1787%now\, \$1705%now\, \$1593_i%now\, \$1853%now\, \$1831_loop99399_result%now\, \$1765_loop99399_arg%now\, \$1710_nb2%now\, \$v581%now\, \$v427%now\, \$1732%now\, \$1585%now\, \$1736%now\, \$1594_id%now\, \$v471%now\, \$1678%now\, \$1592%now\, \$1726_id%now\, \$1697%now\, \$1594_result%now\, \$1850%now\, \$v425%now\, \$1603%now\, \$1681%now\, \$1725_i%now\, \result568%now\, \$1672%now\, \$1790%now\, \$1782%now\, \$1649%now\, \$1623%now\, \$1856%now\, \$1825%now\, \$v539%now\, \$1622%now\, \$v497%now\, \$1583%now\, \$1792_id%now\, \$1751_loop99398_result%now\, \$1751_loop99398_arg%now\, \$1611%now\, \$1734%now\, \$1724%now\, \$v469%now\, \$v470%now\, \$1669%now\, \$1835%now\, \$1693%now\, \$v395%now\, \$v431%now\, \$v559%now\, \$v433%now\, \$v495%now\, \$1673_loop99401_id%now\, \$1691%now\, \$v481%now\, \$1716%now\, \$1601%now\, \$1702%now\, \$v432%now\, \$1625%now\, \$1857_id%now\, \$1745%now\, \$1685_loop99398_id%now\, \$1848%now\, \$1830%now\, \$1742%now\, \result418%now\, \$1692%now\, \$1581%now\, \$1591_x%now\, \$1776_nb2%now\, \$1676%now\, \$v590%now\, \$v478%now\, \$1670%now\, \$1739_loop99401_id%now\, \$1653%now\, \$1699_loop99399_arg%now\, \$1587%now\, \$v516%now\, \$1837%now\, \$v428%now\, \$v473%now\, \$v467%now\, \$1712_loop99400_arg%now\, \$1607_loop99401_id%now\, \$1715%now\, \$v466%now\, \$v562%now\, \$v501%now\, \$v593%now\, \$1659_i%now\, \$1827%now\, \$1617%now\, \$1750_nb2%now\, \$v435%now\, \$1851%now\, \$1743%now\, \$v573%now\, \$1788%now\, \rdy419%now\, \$v520%now\, \$1854%now\, \$v565%now\, \$1805_loop99401_arg%now\, \$1781%now\, \rdy461%now\, \rdy404%now\, \result448%now\, \$v429%now\, \$1694%now\, \$1840%now\, \$1775%now\, \$1629%now\, \$1712_loop99400_result%now\, \$v480%now\, \rdy527%now\, \$v509%now\, \rdy485%now\, \$1778_loop99400_id%now\, \$1588_id%now\, \$1841%now\, \$1817_loop99398_arg%now\, \$v459%now\, \$1792_result%now\, \$1768%now\, \$1632%now\, \$v521%now\, \$v476%now\, \$1598%now\, \$1657_nb2%now\, \$1644_nb2%now\, \$1696_nb2%now\, \$v438%now\, \$v555%now\, \$1718%now\, \$1796%now\, \$1844_loop99400_id%now\, \$v424%now\, \$1584%now\, \$1855_nb2%now\, \$v456%now\, \$1619_loop99398_id%now\, \$1817_loop99398_result%now\, \$1642%now\, \$1619_loop99398_arg%now\, \$v426%now\, \$v397%now\, \$1689%now\, \$1847%now\, \$1679%now\, \result442%now\, \$1844_loop99400_result%now\, \$v537%now\, \$1783%now\, \$v489%now\, \$1809%now\, \$1849%now\, \$1607_loop99401_result%now\, \$v436%now\, \$1826%now\, \$v472%now\, \$v434%now\, \$1602%now\, \$1792_arg%now\, \result407%now\, \$1778_loop99400_result%now\, \$1761%now\, \$1708%now\, \$1599_n%now\, \$v479%now\, \$1748%now\, \$1800%now\, \$1823%now\, \$v554%now\, \$1726_result%now\, \$1626%now\, \$v552%now\, \$1824%now\, \$1695%now\, \$1699_loop99399_id%now\, \$1739_loop99401_result%now\, \$1747%now\, \$v498%now\, \$1650%now\, \$1624%now\, \$1839%now\, \$1651%now\, \$1667%now\, \$1673_loop99401_result%now\, \$1652%now\, \$1646_loop99400_result%now\, \$1802%now\, \$1777%now\, \$1671%now\, \$1757%now\, \$v453%now\, \$1720%now\, \$v563%now\, \$1749%now\, \$v549%now\, \$v585%now\, \$v423%now\, \$1805_loop99401_id%now\, \$1699_loop99399_result%now\, \$1842_nb2%now\, \$1774%now\, \$1723_nb2%now\, \$1633_loop99399_id%now\, \$1612%now\, \$1829%now\, \$1785%now\, \$1733%now\, \$1773%now\, \$v515%now\, \$v439%now\, \$v551%now\, \$1688%now\, \$1582%now\, \$v430%now\, \rdy545%now\, \$1822%now\, \$1654%now\, \$1786%now\, \$1828_nb2%now\, \$1798%now\, \$1778_loop99400_arg%now\, \$1857_result%now\, \$1660_arg%now\, \$1641%now\, \$1769%now\, \rdy449%now\, \$1857_arg%now\, \$1726_arg%now\, \$1610%now\, \$1804%now\, \$1754%now\, \$1759%now\, \$v465%now\, \$v531%now\, \$v508%now\, \$1643%now\, \result490%now\, \$v564%now\, \$1656%now\, \$v437%now\, \$1586%now\, \$1760%now\, \$1813%now\, \$1721%now\, \$1680%now\, \$v522%now\, \$1668%now\, \$1831_loop99399_id%now\, \result526%now\, \$1746%now\, \$v560%now\, \rdy443%now\, \$v475%now\, \$1588_result%now\, \$v477%now\, \$1607_loop99401_arg%now\, \$1631%now\, \$v582%now\, \$v514%now\, \$1772%now\, \$1739_loop99401_arg%now\, \$v455%now\, \$1580_led%now\, \$v587%now\, \$1605%now\, \$1820%now\, \$v468%now\, \rdy575%now\, \$1801%now\, \$1660_result%now\, \$v556%now\, \$1861%now\, \$1764%now\, \$1836%now\, \$1838%now\, \$v558%now\, \$1738%now\, \$1630_nb2%now\, \$1579%now\, \$1805_loop99401_result%now\, \$1729_i%now\, \$1751_loop99398_id%now\, \$1722%now\, \$1618_nb2%now\, \$1795_i%now\, \$1758%now\, \$1658%now\, \$v519%now\, \$1784%now\, \$1763%now\, \$1588_arg%now\, \$1616%now\, \$1808%now\, \result532%now\, \$1655%now\, \$v594%now\, \rdy533%now\, \$1765_loop99399_result%now\, \$v523%now\, \$1604%now\, \$1711%now\, \$1663_i%now\, \$1636%now\, \$1799%now\, \$1810%now\, \$1831_loop99399_arg%now\, \$1731_n%now\, \$v474%now\, \$v510%now\, \$1594_arg%now\, \$1615%now\, \$v518%now\, \$1717%now\, \$1706%now\, \$1606%now\, \$1789_nb2%now\, \$1600%now\, \$1770%now\, \$1709%now\, \$1673_loop99401_arg%now\, \$1704%now\, \$1690%now\, \$1619_loop99398_result%now\, \rdy503%now\, \$1812%now\, \$1614%now\, \$v412%now\, \$$1209_src_lock%now\, \$$1216_dst_lock%now\, \$$1217_r_lock%now\)
        variable \$1614\, \$1812\, \$1690\, \$1704\, \$1709\, \$1770\, 
                 \$1706\, \$1717\, \$1615\, \$1810\, \$1636\, \$1655\, 
                 \$1808\, \$1616\, \$1784\, \$1758\, \$1722\, \$1838\, 
                 \$1836\, \$1820\, \$1772\, \$1746\, \$1680\, \$1721\, 
                 \$1813\, \$1760\, \$1656\, \$1643\, \$1759\, \$1754\, 
                 \$1610\, \$1857_arg\, \$1769\, \$1641\, \$1786\, \$1654\, 
                 \$1822\, \$1688\, \$1773\, \$1785\, \$1612\, \$1774\, 
                 \$1749\, \$1720\, \$1757\, \$1652\, \$1651\, \$1839\, 
                 \$1624\, \$1650\, \$1747\, \$1695\, \$1824\, \$1626\, 
                 \$1823\, \$1748\, \$1708\, \$1761\, \$1826\, \$1849\, 
                 \$1809\, \$1783\, \$1679\, \$1847\, \$1689\, \$1642\, 
                 \$1796\, \$1718\, \$1598\, \$1768\, \$1841\, \$1629\, 
                 \$1775\, \$1840\, \$1694\, \$1781\, \$1854\, \$1788\, 
                 \$1743\, \$1851\, \$1617\, \$1827\, \$1715\, \$1837\, 
                 \$1653\, \$1676\, \$1692\, \$1742\, \$1848\, \$1745\, 
                 \$1625\, \$1702\, \$1716\, \$1691\, \$1693\, \$1835\, 
                 \$1611\, \$1622\, \$1825\, \$1623\, \$1649\, \$1782\, 
                 \$1681\, \$1850\, \$1678\, \$1853\, \$1705\, \$1787\, 
                 \$1852\, \$1639\, \$1628\, \$1771\, \$1815\, \$1638\, 
                 \$1677\, \$1755\, \$1814\, \$1707\, \$1578\, \$1613\, 
                 \$1627\, \$1640\, \$1821\, \$1703\, \$1811\, \$1719\, 
                 \$1756\, \$1730\, \$1637\, \$1683\, \$1834\, \$1682\, 
                 \$1744\, \$1664\ : value(0 to 32) := (others => '0');
        variable \$1594_arg\, \$1726_arg\, \$1660_arg\, \$1792_arg\, \$1592\ : value(0 to 3) := (others => '0');
        variable result403 : value(0 to 57) := (others => '0');
        variable \$1751_loop99398_id\, \$1831_loop99399_id\, 
                 \$1633_loop99399_id\, \$1805_loop99401_id\, 
                 \$1699_loop99399_id\, \$1619_loop99398_id\, 
                 \$1844_loop99400_id\, \$1588_id\, \$1778_loop99400_id\, 
                 \$1607_loop99401_id\, \$1739_loop99401_id\, 
                 \$1685_loop99398_id\, \$1857_id\, \$1673_loop99401_id\, 
                 \$1792_id\, \$1726_id\, \$1594_id\, \$1817_loop99398_id\, 
                 \$1660_id\, \$1712_loop99400_id\, \$1765_loop99399_id\, 
                 \$1646_loop99400_id\ : value(0 to 11) := (others => '0');
        variable \$1588_arg\ : value(0 to 64) := (others => '0');
        variable \$1861\, \$1577_o\ : value(0 to 127) := (others => '0');
        variable \$v412\, rdy503, \$1600\, \$1606\, \$v518\, \$v510\, 
                 \$v474\, \$1799\, \$1711\, \$v523\, rdy533, \$v594\, 
                 \$1763\, \$v519\, \$1658\, \$1579\, \$1738\, \$v558\, 
                 \$1764\, \$v556\, \$1660_result\, \$1801\, rdy575, \$v468\, 
                 \$1605\, \$v587\, \$1580_led\, \$v455\, \$v514\, \$v582\, 
                 \$1631\, \$v477\, \$v475\, rdy443, \$v560\, result526, 
                 \$1668\, \$v522\, \$1586\, \$v437\, \$v564\, \$v508\, 
                 \$v531\, \$v465\, \$1804\, rdy449, \$1857_result\, \$1798\, 
                 rdy545, \$v430\, \$1582\, \$v551\, \$v439\, \$v515\, 
                 \$1733\, \$1829\, \$v423\, \$v585\, \$v549\, \$v563\, 
                 \$v453\, \$1671\, \$1777\, \$1667\, \$v498\, \$v552\, 
                 \$1726_result\, \$v554\, \$1800\, \$v479\, \$1602\, \$v434\, 
                 \$v472\, \$v436\, \$v489\, \$v537\, result442, \$v397\, 
                 \$v426\, \$v456\, \$1584\, \$v424\, \$v555\, \$v438\, 
                 \$v476\, \$v521\, \$1632\, \$1792_result\, \$v459\, rdy485, 
                 \$v509\, rdy527, \$v480\, \$v429\, rdy404, rdy461, \$v565\, 
                 \$v520\, rdy419, \$v573\, \$v435\, \$v593\, \$v501\, 
                 \$v562\, \$v466\, \$v467\, \$v473\, \$v428\, \$v516\, 
                 \$1587\, \$v478\, \$v590\, \$1581\, result418, \$1830\, 
                 \$v432\, \$1601\, \$v481\, \$v495\, \$v433\, \$v559\, 
                 \$v431\, \$v395\, \$1669\, \$v470\, \$v469\, \$1724\, 
                 \$1734\, \$1583\, \$v497\, \$v539\, \$1856\, \$1790\, 
                 \$1672\, result568, \$1603\, \$v425\, \$1594_result\, 
                 \$1697\, \$v471\, \$1585\, \$1732\, \$v427\, \$v581\, 
                 \$1860\, rdy408, rdy491, \$v543\, \$v517\, \$v540\, \$v513\, 
                 result484, \$1843\, \$v406\, \$v507\, result544, \$v550\, 
                 result502, \$v512\, result460, \$1645\, \$v553\, \$v413\, 
                 \$v557\, \$v579\, \$v561\, \$1735\, \$1698\, \$1803\, 
                 \$1666\, \$v447\, \$v596\, \$v511\, \$1737\, rdy569 : value(0 to 0) := (others => '0');
        variable \$1619_loop99398_result\, \$1789_nb2\, \$1731_n\, \$1663_i\, 
                 \$1604\, \$1765_loop99399_result\, result532, \$1795_i\, 
                 \$1618_nb2\, \$1729_i\, \$1805_loop99401_result\, 
                 \$1630_nb2\, \$1588_result\, result490, \$1828_nb2\, 
                 \$1723_nb2\, \$1842_nb2\, \$1699_loop99399_result\, \$1802\, 
                 \$1646_loop99400_result\, \$1673_loop99401_result\, 
                 \$1739_loop99401_result\, \$1599_n\, 
                 \$1778_loop99400_result\, result407, 
                 \$1607_loop99401_result\, \$1844_loop99400_result\, 
                 \$1817_loop99398_result\, \$1855_nb2\, \$1696_nb2\, 
                 \$1644_nb2\, \$1657_nb2\, \$1712_loop99400_result\, 
                 result448, \$1750_nb2\, \$1659_i\, \$1670\, \$1776_nb2\, 
                 \$1591_x\, \$1751_loop99398_result\, \$1725_i\, \$1736\, 
                 \$1710_nb2\, \$1831_loop99399_result\, \$1593_i\, \$1597_i\, 
                 \$1665_n\, \$1791_i\, \$1816_nb2\, \$1684_nb2\, result574, 
                 \$1685_loop99398_result\, \$1797_n\, 
                 \$1633_loop99399_result\, \$1762_nb2\ : value(0 to 31) := (others => '0');
        variable \$1673_loop99401_arg\, \$1831_loop99399_arg\, 
                 \$1739_loop99401_arg\, \$1607_loop99401_arg\, 
                 \$1778_loop99400_arg\, \$1619_loop99398_arg\, 
                 \$1817_loop99398_arg\, \$1805_loop99401_arg\, 
                 \$1712_loop99400_arg\, \$1699_loop99399_arg\, 
                 \$1751_loop99398_arg\, \$1765_loop99399_arg\, 
                 \$1844_loop99400_arg\, \$1633_loop99399_arg\, 
                 \$1646_loop99400_arg\, \$1685_loop99398_arg\ : value(0 to 415) := (others => '0');
        variable state : t_state;
        variable state_var609 : t_state_var609;
        variable state_var608 : t_state_var608;
        variable state_var607 : t_state_var607;
        variable state_var606 : t_state_var606;
        variable state_var605 : t_state_var605;
        variable state_var604 : t_state_var604;
        variable state_var603 : t_state_var603;
        variable state_var602 : t_state_var602;
        variable state_var601 : t_state_var601;
        variable state_var600 : t_state_var600;
        variable state_var599 : t_state_var599;
        variable state_var598 : t_state_var598;
        variable state_var597 : t_state_var597;
        variable \$$1209_src_lock\ : value(0 to 0);
        variable \$$1216_dst_lock\ : value(0 to 0);
        variable \$$1217_r_lock\ : value(0 to 0);
        
    begin
      rdy569 := \rdy569%now\;
      \$1737\ := \$1737%now\;
      \$1646_loop99400_id\ := \$1646_loop99400_id%now\;
      \$1685_loop99398_arg\ := \$1685_loop99398_arg%now\;
      \$v511\ := \$v511%now\;
      \$1664\ := \$1664%now\;
      \$1744\ := \$1744%now\;
      \$1682\ := \$1682%now\;
      \$1762_nb2\ := \$1762_nb2%now\;
      \$v596\ := \$v596%now\;
      \$1577_o\ := \$1577_o%now\;
      \$v447\ := \$v447%now\;
      \$1666\ := \$1666%now\;
      \$1834\ := \$1834%now\;
      \$1683\ := \$1683%now\;
      \$1633_loop99399_result\ := \$1633_loop99399_result%now\;
      \$1637\ := \$1637%now\;
      \$1646_loop99400_arg\ := \$1646_loop99400_arg%now\;
      \$1803\ := \$1803%now\;
      \$1797_n\ := \$1797_n%now\;
      \$1698\ := \$1698%now\;
      \$1735\ := \$1735%now\;
      \$1730\ := \$1730%now\;
      \$1685_loop99398_result\ := \$1685_loop99398_result%now\;
      \$v561\ := \$v561%now\;
      \$1756\ := \$1756%now\;
      \$1765_loop99399_id\ := \$1765_loop99399_id%now\;
      \$v579\ := \$v579%now\;
      \$v557\ := \$v557%now\;
      \$1719\ := \$1719%now\;
      \$v413\ := \$v413%now\;
      \$1811\ := \$1811%now\;
      \$1703\ := \$1703%now\;
      \$1821\ := \$1821%now\;
      \$1640\ := \$1640%now\;
      \$1633_loop99399_arg\ := \$1633_loop99399_arg%now\;
      \$v553\ := \$v553%now\;
      \$1645\ := \$1645%now\;
      \$1627\ := \$1627%now\;
      \$1613\ := \$1613%now\;
      \$1712_loop99400_id\ := \$1712_loop99400_id%now\;
      \$1578\ := \$1578%now\;
      \$1707\ := \$1707%now\;
      \$1814\ := \$1814%now\;
      result574 := \result574%now\;
      \$1755\ := \$1755%now\;
      \$1677\ := \$1677%now\;
      result460 := \result460%now\;
      \$1638\ := \$1638%now\;
      \$v512\ := \$v512%now\;
      result502 := \result502%now\;
      \$1815\ := \$1815%now\;
      \$1771\ := \$1771%now\;
      \$1684_nb2\ := \$1684_nb2%now\;
      \$1660_id\ := \$1660_id%now\;
      \$v550\ := \$v550%now\;
      result544 := \result544%now\;
      \$v507\ := \$v507%now\;
      \$v406\ := \$v406%now\;
      \$1844_loop99400_arg\ := \$1844_loop99400_arg%now\;
      \$1816_nb2\ := \$1816_nb2%now\;
      \$1791_i\ := \$1791_i%now\;
      \$1843\ := \$1843%now\;
      \$1817_loop99398_id\ := \$1817_loop99398_id%now\;
      result484 := \result484%now\;
      \$1628\ := \$1628%now\;
      result403 := \result403%now\;
      \$v513\ := \$v513%now\;
      \$1639\ := \$1639%now\;
      \$v540\ := \$v540%now\;
      \$v517\ := \$v517%now\;
      \$1665_n\ := \$1665_n%now\;
      \$v543\ := \$v543%now\;
      rdy491 := \rdy491%now\;
      rdy408 := \rdy408%now\;
      \$1597_i\ := \$1597_i%now\;
      \$1860\ := \$1860%now\;
      \$1852\ := \$1852%now\;
      \$1787\ := \$1787%now\;
      \$1705\ := \$1705%now\;
      \$1593_i\ := \$1593_i%now\;
      \$1853\ := \$1853%now\;
      \$1831_loop99399_result\ := \$1831_loop99399_result%now\;
      \$1765_loop99399_arg\ := \$1765_loop99399_arg%now\;
      \$1710_nb2\ := \$1710_nb2%now\;
      \$v581\ := \$v581%now\;
      \$v427\ := \$v427%now\;
      \$1732\ := \$1732%now\;
      \$1585\ := \$1585%now\;
      \$1736\ := \$1736%now\;
      \$1594_id\ := \$1594_id%now\;
      \$v471\ := \$v471%now\;
      \$1678\ := \$1678%now\;
      \$1592\ := \$1592%now\;
      \$1726_id\ := \$1726_id%now\;
      \$1697\ := \$1697%now\;
      \$1594_result\ := \$1594_result%now\;
      \$1850\ := \$1850%now\;
      \$v425\ := \$v425%now\;
      \$1603\ := \$1603%now\;
      \$1681\ := \$1681%now\;
      \$1725_i\ := \$1725_i%now\;
      result568 := \result568%now\;
      \$1672\ := \$1672%now\;
      \$1790\ := \$1790%now\;
      \$1782\ := \$1782%now\;
      \$1649\ := \$1649%now\;
      \$1623\ := \$1623%now\;
      \$1856\ := \$1856%now\;
      \$1825\ := \$1825%now\;
      \$v539\ := \$v539%now\;
      \$1622\ := \$1622%now\;
      \$v497\ := \$v497%now\;
      \$1583\ := \$1583%now\;
      \$1792_id\ := \$1792_id%now\;
      \$1751_loop99398_result\ := \$1751_loop99398_result%now\;
      \$1751_loop99398_arg\ := \$1751_loop99398_arg%now\;
      \$1611\ := \$1611%now\;
      \$1734\ := \$1734%now\;
      \$1724\ := \$1724%now\;
      \$v469\ := \$v469%now\;
      \$v470\ := \$v470%now\;
      \$1669\ := \$1669%now\;
      \$1835\ := \$1835%now\;
      \$1693\ := \$1693%now\;
      \$v395\ := \$v395%now\;
      \$v431\ := \$v431%now\;
      \$v559\ := \$v559%now\;
      \$v433\ := \$v433%now\;
      \$v495\ := \$v495%now\;
      \$1673_loop99401_id\ := \$1673_loop99401_id%now\;
      \$1691\ := \$1691%now\;
      \$v481\ := \$v481%now\;
      \$1716\ := \$1716%now\;
      \$1601\ := \$1601%now\;
      \$1702\ := \$1702%now\;
      \$v432\ := \$v432%now\;
      \$1625\ := \$1625%now\;
      \$1857_id\ := \$1857_id%now\;
      \$1745\ := \$1745%now\;
      \$1685_loop99398_id\ := \$1685_loop99398_id%now\;
      \$1848\ := \$1848%now\;
      \$1830\ := \$1830%now\;
      \$1742\ := \$1742%now\;
      result418 := \result418%now\;
      \$1692\ := \$1692%now\;
      \$1581\ := \$1581%now\;
      \$1591_x\ := \$1591_x%now\;
      \$1776_nb2\ := \$1776_nb2%now\;
      \$1676\ := \$1676%now\;
      \$v590\ := \$v590%now\;
      \$v478\ := \$v478%now\;
      \$1670\ := \$1670%now\;
      \$1739_loop99401_id\ := \$1739_loop99401_id%now\;
      \$1653\ := \$1653%now\;
      \$1699_loop99399_arg\ := \$1699_loop99399_arg%now\;
      \$1587\ := \$1587%now\;
      \$v516\ := \$v516%now\;
      \$1837\ := \$1837%now\;
      \$v428\ := \$v428%now\;
      \$v473\ := \$v473%now\;
      \$v467\ := \$v467%now\;
      \$1712_loop99400_arg\ := \$1712_loop99400_arg%now\;
      \$1607_loop99401_id\ := \$1607_loop99401_id%now\;
      \$1715\ := \$1715%now\;
      \$v466\ := \$v466%now\;
      \$v562\ := \$v562%now\;
      \$v501\ := \$v501%now\;
      \$v593\ := \$v593%now\;
      \$1659_i\ := \$1659_i%now\;
      \$1827\ := \$1827%now\;
      \$1617\ := \$1617%now\;
      \$1750_nb2\ := \$1750_nb2%now\;
      \$v435\ := \$v435%now\;
      \$1851\ := \$1851%now\;
      \$1743\ := \$1743%now\;
      \$v573\ := \$v573%now\;
      \$1788\ := \$1788%now\;
      rdy419 := \rdy419%now\;
      \$v520\ := \$v520%now\;
      \$1854\ := \$1854%now\;
      \$v565\ := \$v565%now\;
      \$1805_loop99401_arg\ := \$1805_loop99401_arg%now\;
      \$1781\ := \$1781%now\;
      rdy461 := \rdy461%now\;
      rdy404 := \rdy404%now\;
      result448 := \result448%now\;
      \$v429\ := \$v429%now\;
      \$1694\ := \$1694%now\;
      \$1840\ := \$1840%now\;
      \$1775\ := \$1775%now\;
      \$1629\ := \$1629%now\;
      \$1712_loop99400_result\ := \$1712_loop99400_result%now\;
      \$v480\ := \$v480%now\;
      rdy527 := \rdy527%now\;
      \$v509\ := \$v509%now\;
      rdy485 := \rdy485%now\;
      \$1778_loop99400_id\ := \$1778_loop99400_id%now\;
      \$1588_id\ := \$1588_id%now\;
      \$1841\ := \$1841%now\;
      \$1817_loop99398_arg\ := \$1817_loop99398_arg%now\;
      \$v459\ := \$v459%now\;
      \$1792_result\ := \$1792_result%now\;
      \$1768\ := \$1768%now\;
      \$1632\ := \$1632%now\;
      \$v521\ := \$v521%now\;
      \$v476\ := \$v476%now\;
      \$1598\ := \$1598%now\;
      \$1657_nb2\ := \$1657_nb2%now\;
      \$1644_nb2\ := \$1644_nb2%now\;
      \$1696_nb2\ := \$1696_nb2%now\;
      \$v438\ := \$v438%now\;
      \$v555\ := \$v555%now\;
      \$1718\ := \$1718%now\;
      \$1796\ := \$1796%now\;
      \$1844_loop99400_id\ := \$1844_loop99400_id%now\;
      \$v424\ := \$v424%now\;
      \$1584\ := \$1584%now\;
      \$1855_nb2\ := \$1855_nb2%now\;
      \$v456\ := \$v456%now\;
      \$1619_loop99398_id\ := \$1619_loop99398_id%now\;
      \$1817_loop99398_result\ := \$1817_loop99398_result%now\;
      \$1642\ := \$1642%now\;
      \$1619_loop99398_arg\ := \$1619_loop99398_arg%now\;
      \$v426\ := \$v426%now\;
      \$v397\ := \$v397%now\;
      \$1689\ := \$1689%now\;
      \$1847\ := \$1847%now\;
      \$1679\ := \$1679%now\;
      result442 := \result442%now\;
      \$1844_loop99400_result\ := \$1844_loop99400_result%now\;
      \$v537\ := \$v537%now\;
      \$1783\ := \$1783%now\;
      \$v489\ := \$v489%now\;
      \$1809\ := \$1809%now\;
      \$1849\ := \$1849%now\;
      \$1607_loop99401_result\ := \$1607_loop99401_result%now\;
      \$v436\ := \$v436%now\;
      \$1826\ := \$1826%now\;
      \$v472\ := \$v472%now\;
      \$v434\ := \$v434%now\;
      \$1602\ := \$1602%now\;
      \$1792_arg\ := \$1792_arg%now\;
      result407 := \result407%now\;
      \$1778_loop99400_result\ := \$1778_loop99400_result%now\;
      \$1761\ := \$1761%now\;
      \$1708\ := \$1708%now\;
      \$1599_n\ := \$1599_n%now\;
      \$v479\ := \$v479%now\;
      \$1748\ := \$1748%now\;
      \$1800\ := \$1800%now\;
      \$1823\ := \$1823%now\;
      \$v554\ := \$v554%now\;
      \$1726_result\ := \$1726_result%now\;
      \$1626\ := \$1626%now\;
      \$v552\ := \$v552%now\;
      \$1824\ := \$1824%now\;
      \$1695\ := \$1695%now\;
      \$1699_loop99399_id\ := \$1699_loop99399_id%now\;
      \$1739_loop99401_result\ := \$1739_loop99401_result%now\;
      \$1747\ := \$1747%now\;
      \$v498\ := \$v498%now\;
      \$1650\ := \$1650%now\;
      \$1624\ := \$1624%now\;
      \$1839\ := \$1839%now\;
      \$1651\ := \$1651%now\;
      \$1667\ := \$1667%now\;
      \$1673_loop99401_result\ := \$1673_loop99401_result%now\;
      \$1652\ := \$1652%now\;
      \$1646_loop99400_result\ := \$1646_loop99400_result%now\;
      \$1802\ := \$1802%now\;
      \$1777\ := \$1777%now\;
      \$1671\ := \$1671%now\;
      \$1757\ := \$1757%now\;
      \$v453\ := \$v453%now\;
      \$1720\ := \$1720%now\;
      \$v563\ := \$v563%now\;
      \$1749\ := \$1749%now\;
      \$v549\ := \$v549%now\;
      \$v585\ := \$v585%now\;
      \$v423\ := \$v423%now\;
      \$1805_loop99401_id\ := \$1805_loop99401_id%now\;
      \$1699_loop99399_result\ := \$1699_loop99399_result%now\;
      \$1842_nb2\ := \$1842_nb2%now\;
      \$1774\ := \$1774%now\;
      \$1723_nb2\ := \$1723_nb2%now\;
      \$1633_loop99399_id\ := \$1633_loop99399_id%now\;
      \$1612\ := \$1612%now\;
      \$1829\ := \$1829%now\;
      \$1785\ := \$1785%now\;
      \$1733\ := \$1733%now\;
      \$1773\ := \$1773%now\;
      \$v515\ := \$v515%now\;
      \$v439\ := \$v439%now\;
      \$v551\ := \$v551%now\;
      \$1688\ := \$1688%now\;
      \$1582\ := \$1582%now\;
      \$v430\ := \$v430%now\;
      rdy545 := \rdy545%now\;
      \$1822\ := \$1822%now\;
      \$1654\ := \$1654%now\;
      \$1786\ := \$1786%now\;
      \$1828_nb2\ := \$1828_nb2%now\;
      \$1798\ := \$1798%now\;
      \$1778_loop99400_arg\ := \$1778_loop99400_arg%now\;
      \$1857_result\ := \$1857_result%now\;
      \$1660_arg\ := \$1660_arg%now\;
      \$1641\ := \$1641%now\;
      \$1769\ := \$1769%now\;
      rdy449 := \rdy449%now\;
      \$1857_arg\ := \$1857_arg%now\;
      \$1726_arg\ := \$1726_arg%now\;
      \$1610\ := \$1610%now\;
      \$1804\ := \$1804%now\;
      \$1754\ := \$1754%now\;
      \$1759\ := \$1759%now\;
      \$v465\ := \$v465%now\;
      \$v531\ := \$v531%now\;
      \$v508\ := \$v508%now\;
      \$1643\ := \$1643%now\;
      result490 := \result490%now\;
      \$v564\ := \$v564%now\;
      \$1656\ := \$1656%now\;
      \$v437\ := \$v437%now\;
      \$1586\ := \$1586%now\;
      \$1760\ := \$1760%now\;
      \$1813\ := \$1813%now\;
      \$1721\ := \$1721%now\;
      \$1680\ := \$1680%now\;
      \$v522\ := \$v522%now\;
      \$1668\ := \$1668%now\;
      \$1831_loop99399_id\ := \$1831_loop99399_id%now\;
      result526 := \result526%now\;
      \$1746\ := \$1746%now\;
      \$v560\ := \$v560%now\;
      rdy443 := \rdy443%now\;
      \$v475\ := \$v475%now\;
      \$1588_result\ := \$1588_result%now\;
      \$v477\ := \$v477%now\;
      \$1607_loop99401_arg\ := \$1607_loop99401_arg%now\;
      \$1631\ := \$1631%now\;
      \$v582\ := \$v582%now\;
      \$v514\ := \$v514%now\;
      \$1772\ := \$1772%now\;
      \$1739_loop99401_arg\ := \$1739_loop99401_arg%now\;
      \$v455\ := \$v455%now\;
      \$1580_led\ := \$1580_led%now\;
      \$v587\ := \$v587%now\;
      \$1605\ := \$1605%now\;
      \$1820\ := \$1820%now\;
      \$v468\ := \$v468%now\;
      rdy575 := \rdy575%now\;
      \$1801\ := \$1801%now\;
      \$1660_result\ := \$1660_result%now\;
      \$v556\ := \$v556%now\;
      \$1861\ := \$1861%now\;
      \$1764\ := \$1764%now\;
      \$1836\ := \$1836%now\;
      \$1838\ := \$1838%now\;
      \$v558\ := \$v558%now\;
      \$1738\ := \$1738%now\;
      \$1630_nb2\ := \$1630_nb2%now\;
      \$1579\ := \$1579%now\;
      \$1805_loop99401_result\ := \$1805_loop99401_result%now\;
      \$1729_i\ := \$1729_i%now\;
      \$1751_loop99398_id\ := \$1751_loop99398_id%now\;
      \$1722\ := \$1722%now\;
      \$1618_nb2\ := \$1618_nb2%now\;
      \$1795_i\ := \$1795_i%now\;
      \$1758\ := \$1758%now\;
      \$1658\ := \$1658%now\;
      \$v519\ := \$v519%now\;
      \$1784\ := \$1784%now\;
      \$1763\ := \$1763%now\;
      \$1588_arg\ := \$1588_arg%now\;
      \$1616\ := \$1616%now\;
      \$1808\ := \$1808%now\;
      result532 := \result532%now\;
      \$1655\ := \$1655%now\;
      \$v594\ := \$v594%now\;
      rdy533 := \rdy533%now\;
      \$1765_loop99399_result\ := \$1765_loop99399_result%now\;
      \$v523\ := \$v523%now\;
      \$1604\ := \$1604%now\;
      \$1711\ := \$1711%now\;
      \$1663_i\ := \$1663_i%now\;
      \$1636\ := \$1636%now\;
      \$1799\ := \$1799%now\;
      \$1810\ := \$1810%now\;
      \$1831_loop99399_arg\ := \$1831_loop99399_arg%now\;
      \$1731_n\ := \$1731_n%now\;
      \$v474\ := \$v474%now\;
      \$v510\ := \$v510%now\;
      \$1594_arg\ := \$1594_arg%now\;
      \$1615\ := \$1615%now\;
      \$v518\ := \$v518%now\;
      \$1717\ := \$1717%now\;
      \$1706\ := \$1706%now\;
      \$1606\ := \$1606%now\;
      \$1789_nb2\ := \$1789_nb2%now\;
      \$1600\ := \$1600%now\;
      \$1770\ := \$1770%now\;
      \$1709\ := \$1709%now\;
      \$1673_loop99401_arg\ := \$1673_loop99401_arg%now\;
      \$1704\ := \$1704%now\;
      \$1690\ := \$1690%now\;
      \$1619_loop99398_result\ := \$1619_loop99398_result%now\;
      rdy503 := \rdy503%now\;
      \$1812\ := \$1812%now\;
      \$1614\ := \$1614%now\;
      \$v412\ := \$v412%now\;
      \$$1209_src_lock\ := \$$1209_src_lock%now\;
      \$$1216_dst_lock\ := \$$1216_dst_lock%now\;
      \$$1217_r_lock\ := \$$1217_r_lock%now\;
      state := \state%now\;
      state_var609 := \state_var609%now\;
      state_var608 := \state_var608%now\;
      state_var607 := \state_var607%now\;
      state_var606 := \state_var606%now\;
      state_var605 := \state_var605%now\;
      state_var604 := \state_var604%now\;
      state_var603 := \state_var603%now\;
      state_var602 := \state_var602%now\;
      state_var601 := \state_var601%now\;
      state_var600 := \state_var600%now\;
      state_var599 := \state_var599%now\;
      state_var598 := \state_var598%now\;
      state_var597 := \state_var597%now\;
      case state is
      when IDLE405 =>
        rdy404 := eclat_false;
        \$v596\ := eclat_if(""&argument(0) & eclat_true & ""&argument(1));
        if \$v596\(0) = '1' then
          result403 := eclat_true & "0"& X"0000000000000" & X"0";
          rdy404 := eclat_true;
          state := IDLE405;
        else
          if \$v395\(0) = '1' then
            
          else
            \$v395\ := eclat_true;
            \$1861\ := work.Int.neg(X"0000000000000000000000000000000" & X"1");
          end if;
          \$1861\ := work.Int.add(\$1861\, X"0000000000000000000000000000000" & X"1");
          \$1577_o\ := \$1861\;
          case state_var597 is
          when \$1588\ =>
            \$v413\ := work.Int.lt(\$1588_arg\(32 to 63), std_logic_vector(to_unsigned(\$1216_dst\'length,32)));
            if \$v413\(0) = '1' then
              \$v412\ := \$$1216_dst_lock\;
              if \$v412\(0) = '1' then
                state_var597 := Q_WAIT411;
              else
                acquire(\$$1216_dst_lock\);
                \$$1216_dst_ptr\ <= to_integer(unsigned(\$1588_arg\(32 to 63)));
                state_var597 := PAUSE_GET410;
              end if;
            else
              \$1588_result\ := \$1588_arg\(0 to 31);
              result407 := \$1588_result\;
              rdy408 := eclat_true;
              state_var597 := IDLE409;
            end if;
          when \$1857\ =>
            \$v594\ := work.Int.gt(\$1857_arg\(0 to 31), work.Int.sub(
                                                         std_logic_vector(to_unsigned(\$1209_src\'length,32)), X"0000000" & X"1"));
            if \$v594\(0) = '1' then
              \$1857_result\ := eclat_unit;
              \$1585\ := \$1857_result\;
              \$v590\ := \$$1217_r_lock\;
              if \$v590\(0) = '1' then
                state_var597 := Q_WAIT589;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= X"0000000" & X"0"; \$$1217_r_write_request\ <= '1';
                state_var597 := PAUSE_SET588;
              end if;
            else
              \$v593\ := \$$1209_src_lock\;
              if \$v593\(0) = '1' then
                state_var597 := Q_WAIT592;
              else
                acquire(\$$1209_src_lock\);
                \$$1209_src_ptr_write\ <= to_integer(unsigned(\$1857_arg\(0 to 31)));
                \$$1209_src_write\ <= work.Int.add(\$1857_arg\(0 to 31), X"0000000" & X"1"); \$$1209_src_write_request\ <= '1';
                state_var597 := PAUSE_SET591;
              end if;
            end if;
          when PAR586 =>
            case state_var607 is
            when \$1594\ =>
              \$v459\ := \$$1217_r_lock\;
              if \$v459\(0) = '1' then
                state_var607 := Q_WAIT458;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var607 := PAUSE_GET457;
              end if;
            when \$1607_LOOP99401\ =>
              \$v439\ := work.Int.le(\$1607_loop99401_arg\(64 to 95), \$1607_loop99401_arg\(96 to 127));
              if \$v439\(0) = '1' then
                \$1617\ := X"0000000" & X"7" & eclat_true;
                \$1616\ := X"0000000" & X"6" & work.Bool.land(""&\$1617\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1617\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1617\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1617\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1617\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1617\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1617\(0 to 31))) & eclat_false)));
                \$1615\ := X"0000000" & X"5" & work.Bool.land(""&\$1616\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1616\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1616\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1616\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1616\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1616\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1616\(0 to 31))) & eclat_false)));
                \$1614\ := X"0000000" & X"4" & work.Bool.land(""&\$1615\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1615\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1615\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1615\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1615\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1615\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1615\(0 to 31))) & eclat_false)));
                \$1613\ := X"0000000" & X"3" & work.Bool.land(""&\$1614\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1614\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1614\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1614\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1614\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1614\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1614\(0 to 31))) & eclat_false)));
                \$1612\ := X"0000000" & X"2" & work.Bool.land(""&\$1613\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1613\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1613\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1613\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1613\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1613\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1613\(0 to 31))) & eclat_false)));
                \$1611\ := X"0000000" & X"1" & work.Bool.land(""&\$1612\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1612\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1612\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1612\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1612\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1612\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1612\(0 to 31))) & eclat_false)));
                \$1610\ := X"0000000" & X"0" & work.Bool.land(""&\$1611\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1611\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1611\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1611\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1611\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1611\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1607_loop99401_arg\(32 to 63), \$1611\(0 to 31))) & eclat_false)));
                \$v433\ := work.Bool.land(""&\$1610\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1610\(0 to 31), X"0000000" & X"1"), \$1607_loop99401_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1610\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1610\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1610\(0 to 31),16),16)), \$1607_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1607_loop99401_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1610\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1607_loop99401_arg\(32 to 63), \$1610\(0 to 31))) & eclat_false)));
                if \$v433\(0) = '1' then
                  \$v428\ := work.Int.eq(work.Int.add(\$1607_loop99401_arg\(32 to 63), X"0000000" & X"1"), \$1607_loop99401_arg\(96 to 127));
                  if \$v428\(0) = '1' then
                    \$1632\ := work.Print.print_string(clk,of_string("foo"));
                    \$1618_nb2\ := work.Int.add(\$1607_loop99401_arg\(384 to 415), X"0000000" & X"1");
                    \$1619_loop99398_id\ := "000000000010";
                    \$1619_loop99398_arg\ := \$1607_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1607_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1607_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1607_loop99401_arg\(32 to 63),32),16), \$1607_loop99401_arg\(64 to 95)) & \$1618_nb2\;
                    state_var607 := \$1619_LOOP99398\;
                  else
                    \$1618_nb2\ := \$1607_loop99401_arg\(384 to 415);
                    \$1619_loop99398_id\ := "000000000010";
                    \$1619_loop99398_arg\ := \$1607_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1607_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1607_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1607_loop99401_arg\(32 to 63),32),16), \$1607_loop99401_arg\(64 to 95)) & \$1618_nb2\;
                    state_var607 := \$1619_LOOP99398\;
                  end if;
                else
                  \$1633_loop99399_id\ := "000000000011";
                  \$1633_loop99399_arg\ := \$1607_loop99401_arg\(0 to 31) & \$1607_loop99401_arg\(32 to 63) & 
                  work.Int.add(\$1607_loop99401_arg\(64 to 95), X"0000000" & X"1") & \$1607_loop99401_arg\(96 to 127) & \$1607_loop99401_arg\(128 to 383) & \$1607_loop99401_arg\(384 to 415);
                  state_var607 := \$1633_LOOP99399\;
                end if;
              else
                \$v438\ := work.Int.ge(\$1607_loop99401_arg\(32 to 63), \$1607_loop99401_arg\(0 to 31));
                if \$v438\(0) = '1' then
                  \$1646_loop99400_id\ := "000000000100";
                  \$1646_loop99400_arg\ := \$1607_loop99401_arg\(0 to 31) & 
                  work.Int.sub(\$1607_loop99401_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1607_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1607_loop99401_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1607_loop99401_arg\(96 to 127) & \$1607_loop99401_arg\(128 to 383) & \$1607_loop99401_arg\(384 to 415);
                  state_var607 := \$1646_LOOP99400\;
                else
                  \$1607_loop99401_result\ := \$1607_loop99401_arg\(384 to 415);
                  \$1599_n\ := \$1607_loop99401_result\;
                  \$1600\ := work.Print.print_string(clk,of_string("rang "));
                  \$1601\ := work.Int.print(clk,\$1598\(1 to 32));
                  \$1602\ := work.Print.print_string(clk,of_string(": "));
                  \$1603\ := work.Int.print(clk,\$1599_n\);
                  \$1606\ := work.Print.print_newline(clk,eclat_unit);
                  \$1604\ := \$1599_n\;
                  \$v423\ := \$$1216_dst_lock\;
                  if \$v423\(0) = '1' then
                    state_var607 := Q_WAIT422;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1597_i\));
                    \$$1216_dst_write\ <= \$1604\; \$$1216_dst_write_request\ <= '1';
                    state_var607 := PAUSE_SET421;
                  end if;
                end if;
              end if;
            when \$1619_LOOP99398\ =>
              \$v427\ := work.Int.le(\$1619_loop99398_arg\(64 to 95), \$1619_loop99398_arg\(96 to 127));
              if \$v427\(0) = '1' then
                \$1629\ := X"0000000" & X"7" & eclat_true;
                \$1628\ := X"0000000" & X"6" & work.Bool.land(""&\$1629\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1629\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1629\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1629\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1629\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1629\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1629\(0 to 31))) & eclat_false)));
                \$1627\ := X"0000000" & X"5" & work.Bool.land(""&\$1628\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1628\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1628\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1628\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1628\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1628\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1628\(0 to 31))) & eclat_false)));
                \$1626\ := X"0000000" & X"4" & work.Bool.land(""&\$1627\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1627\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1627\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1627\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1627\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1627\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1627\(0 to 31))) & eclat_false)));
                \$1625\ := X"0000000" & X"3" & work.Bool.land(""&\$1626\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1626\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1626\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1626\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1626\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1626\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1626\(0 to 31))) & eclat_false)));
                \$1624\ := X"0000000" & X"2" & work.Bool.land(""&\$1625\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1625\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1625\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1625\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1625\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1625\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1625\(0 to 31))) & eclat_false)));
                \$1623\ := X"0000000" & X"1" & work.Bool.land(""&\$1624\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1624\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1624\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1624\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1624\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1624\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1624\(0 to 31))) & eclat_false)));
                \$1622\ := X"0000000" & X"0" & work.Bool.land(""&\$1623\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1623\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1623\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1623\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1623\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1623\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1619_loop99398_arg\(32 to 63), \$1623\(0 to 31))) & eclat_false)));
                \$v425\ := work.Bool.land(""&\$1622\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1622\(0 to 31), X"0000000" & X"1"), \$1619_loop99398_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1622\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1622\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1622\(0 to 31),16),16)), \$1619_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1619_loop99398_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1622\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1619_loop99398_arg\(32 to 63), \$1622\(0 to 31))) & eclat_false)));
                if \$v425\(0) = '1' then
                  \$v424\ := work.Int.eq(work.Int.add(\$1619_loop99398_arg\(32 to 63), X"0000000" & X"1"), \$1619_loop99398_arg\(96 to 127));
                  if \$v424\(0) = '1' then
                    \$1631\ := work.Print.print_string(clk,of_string("foo"));
                    \$1630_nb2\ := work.Int.add(\$1619_loop99398_arg\(384 to 415), X"0000000" & X"1");
                    \$1619_loop99398_arg\ := \$1619_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1619_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1619_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1619_loop99398_arg\(32 to 63),32),16), \$1619_loop99398_arg\(64 to 95)) & \$1630_nb2\;
                    state_var607 := \$1619_LOOP99398\;
                  else
                    \$1630_nb2\ := \$1619_loop99398_arg\(384 to 415);
                    \$1619_loop99398_arg\ := \$1619_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1619_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1619_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1619_loop99398_arg\(32 to 63),32),16), \$1619_loop99398_arg\(64 to 95)) & \$1630_nb2\;
                    state_var607 := \$1619_LOOP99398\;
                  end if;
                else
                  \$1619_loop99398_arg\ := \$1619_loop99398_arg\(0 to 31) & \$1619_loop99398_arg\(32 to 63) & 
                  work.Int.add(\$1619_loop99398_arg\(64 to 95), X"0000000" & X"1") & \$1619_loop99398_arg\(96 to 127) & \$1619_loop99398_arg\(128 to 383) & \$1619_loop99398_arg\(384 to 415);
                  state_var607 := \$1619_LOOP99398\;
                end if;
              else
                \$v426\ := work.Int.ge(\$1619_loop99398_arg\(32 to 63), \$1619_loop99398_arg\(0 to 31));
                if \$v426\(0) = '1' then
                  \$1619_loop99398_arg\ := \$1619_loop99398_arg\(0 to 31) & 
                  work.Int.sub(\$1619_loop99398_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1619_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1619_loop99398_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1619_loop99398_arg\(96 to 127) & \$1619_loop99398_arg\(128 to 383) & \$1619_loop99398_arg\(384 to 415);
                  state_var607 := \$1619_LOOP99398\;
                else
                  \$1619_loop99398_result\ := \$1619_loop99398_arg\(384 to 415);
                  \$1607_loop99401_result\ := \$1619_loop99398_result\;
                  \$1599_n\ := \$1607_loop99401_result\;
                  \$1600\ := work.Print.print_string(clk,of_string("rang "));
                  \$1601\ := work.Int.print(clk,\$1598\(1 to 32));
                  \$1602\ := work.Print.print_string(clk,of_string(": "));
                  \$1603\ := work.Int.print(clk,\$1599_n\);
                  \$1606\ := work.Print.print_newline(clk,eclat_unit);
                  \$1604\ := \$1599_n\;
                  \$v423\ := \$$1216_dst_lock\;
                  if \$v423\(0) = '1' then
                    state_var607 := Q_WAIT422;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1597_i\));
                    \$$1216_dst_write\ <= \$1604\; \$$1216_dst_write_request\ <= '1';
                    state_var607 := PAUSE_SET421;
                  end if;
                end if;
              end if;
            when \$1633_LOOP99399\ =>
              \$v432\ := work.Int.le(\$1633_loop99399_arg\(64 to 95), \$1633_loop99399_arg\(96 to 127));
              if \$v432\(0) = '1' then
                \$1643\ := X"0000000" & X"7" & eclat_true;
                \$1642\ := X"0000000" & X"6" & work.Bool.land(""&\$1643\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1643\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1643\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1643\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1643\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1643\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1643\(0 to 31))) & eclat_false)));
                \$1641\ := X"0000000" & X"5" & work.Bool.land(""&\$1642\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1642\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1642\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1642\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1642\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1642\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1642\(0 to 31))) & eclat_false)));
                \$1640\ := X"0000000" & X"4" & work.Bool.land(""&\$1641\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1641\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1641\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1641\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1641\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1641\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1641\(0 to 31))) & eclat_false)));
                \$1639\ := X"0000000" & X"3" & work.Bool.land(""&\$1640\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1640\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1640\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1640\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1640\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1640\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1640\(0 to 31))) & eclat_false)));
                \$1638\ := X"0000000" & X"2" & work.Bool.land(""&\$1639\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1639\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1639\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1639\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1639\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1639\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1639\(0 to 31))) & eclat_false)));
                \$1637\ := X"0000000" & X"1" & work.Bool.land(""&\$1638\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1638\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1638\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1638\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1638\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1638\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1638\(0 to 31))) & eclat_false)));
                \$1636\ := X"0000000" & X"0" & work.Bool.land(""&\$1637\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1637\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1637\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1637\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1637\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1637\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1633_loop99399_arg\(32 to 63), \$1637\(0 to 31))) & eclat_false)));
                \$v430\ := work.Bool.land(""&\$1636\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1636\(0 to 31), X"0000000" & X"1"), \$1633_loop99399_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1636\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1636\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1636\(0 to 31),16),16)), \$1633_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1633_loop99399_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1636\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1633_loop99399_arg\(32 to 63), \$1636\(0 to 31))) & eclat_false)));
                if \$v430\(0) = '1' then
                  \$v429\ := work.Int.eq(work.Int.add(\$1633_loop99399_arg\(32 to 63), X"0000000" & X"1"), \$1633_loop99399_arg\(96 to 127));
                  if \$v429\(0) = '1' then
                    \$1645\ := work.Print.print_string(clk,of_string("foo"));
                    \$1644_nb2\ := work.Int.add(\$1633_loop99399_arg\(384 to 415), X"0000000" & X"1");
                    \$1633_loop99399_arg\ := \$1633_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1633_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1633_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1633_loop99399_arg\(32 to 63),32),16), \$1633_loop99399_arg\(64 to 95)) & \$1644_nb2\;
                    state_var607 := \$1633_LOOP99399\;
                  else
                    \$1644_nb2\ := \$1633_loop99399_arg\(384 to 415);
                    \$1633_loop99399_arg\ := \$1633_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1633_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1633_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1633_loop99399_arg\(32 to 63),32),16), \$1633_loop99399_arg\(64 to 95)) & \$1644_nb2\;
                    state_var607 := \$1633_LOOP99399\;
                  end if;
                else
                  \$1633_loop99399_arg\ := \$1633_loop99399_arg\(0 to 31) & \$1633_loop99399_arg\(32 to 63) & 
                  work.Int.add(\$1633_loop99399_arg\(64 to 95), X"0000000" & X"1") & \$1633_loop99399_arg\(96 to 127) & \$1633_loop99399_arg\(128 to 383) & \$1633_loop99399_arg\(384 to 415);
                  state_var607 := \$1633_LOOP99399\;
                end if;
              else
                \$v431\ := work.Int.ge(\$1633_loop99399_arg\(32 to 63), \$1633_loop99399_arg\(0 to 31));
                if \$v431\(0) = '1' then
                  \$1633_loop99399_arg\ := \$1633_loop99399_arg\(0 to 31) & 
                  work.Int.sub(\$1633_loop99399_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1633_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1633_loop99399_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1633_loop99399_arg\(96 to 127) & \$1633_loop99399_arg\(128 to 383) & \$1633_loop99399_arg\(384 to 415);
                  state_var607 := \$1633_LOOP99399\;
                else
                  \$1633_loop99399_result\ := \$1633_loop99399_arg\(384 to 415);
                  \$1607_loop99401_result\ := \$1633_loop99399_result\;
                  \$1599_n\ := \$1607_loop99401_result\;
                  \$1600\ := work.Print.print_string(clk,of_string("rang "));
                  \$1601\ := work.Int.print(clk,\$1598\(1 to 32));
                  \$1602\ := work.Print.print_string(clk,of_string(": "));
                  \$1603\ := work.Int.print(clk,\$1599_n\);
                  \$1606\ := work.Print.print_newline(clk,eclat_unit);
                  \$1604\ := \$1599_n\;
                  \$v423\ := \$$1216_dst_lock\;
                  if \$v423\(0) = '1' then
                    state_var607 := Q_WAIT422;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1597_i\));
                    \$$1216_dst_write\ <= \$1604\; \$$1216_dst_write_request\ <= '1';
                    state_var607 := PAUSE_SET421;
                  end if;
                end if;
              end if;
            when \$1646_LOOP99400\ =>
              \$v437\ := work.Int.le(\$1646_loop99400_arg\(64 to 95), \$1646_loop99400_arg\(96 to 127));
              if \$v437\(0) = '1' then
                \$1656\ := X"0000000" & X"7" & eclat_true;
                \$1655\ := X"0000000" & X"6" & work.Bool.land(""&\$1656\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1656\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1656\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1656\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1656\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1656\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1656\(0 to 31))) & eclat_false)));
                \$1654\ := X"0000000" & X"5" & work.Bool.land(""&\$1655\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1655\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1655\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1655\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1655\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1655\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1655\(0 to 31))) & eclat_false)));
                \$1653\ := X"0000000" & X"4" & work.Bool.land(""&\$1654\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1654\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1654\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1654\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1654\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1654\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1654\(0 to 31))) & eclat_false)));
                \$1652\ := X"0000000" & X"3" & work.Bool.land(""&\$1653\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1653\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1653\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1653\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1653\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1653\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1653\(0 to 31))) & eclat_false)));
                \$1651\ := X"0000000" & X"2" & work.Bool.land(""&\$1652\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1652\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1652\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1652\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1652\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1652\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1652\(0 to 31))) & eclat_false)));
                \$1650\ := X"0000000" & X"1" & work.Bool.land(""&\$1651\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1651\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1651\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1651\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1651\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1651\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1651\(0 to 31))) & eclat_false)));
                \$1649\ := X"0000000" & X"0" & work.Bool.land(""&\$1650\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1650\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1650\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1650\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1650\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1650\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1646_loop99400_arg\(32 to 63), \$1650\(0 to 31))) & eclat_false)));
                \$v435\ := work.Bool.land(""&\$1649\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1649\(0 to 31), X"0000000" & X"1"), \$1646_loop99400_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1649\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1649\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1649\(0 to 31),16),16)), \$1646_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1646_loop99400_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1649\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1646_loop99400_arg\(32 to 63), \$1649\(0 to 31))) & eclat_false)));
                if \$v435\(0) = '1' then
                  \$v434\ := work.Int.eq(work.Int.add(\$1646_loop99400_arg\(32 to 63), X"0000000" & X"1"), \$1646_loop99400_arg\(96 to 127));
                  if \$v434\(0) = '1' then
                    \$1658\ := work.Print.print_string(clk,of_string("foo"));
                    \$1657_nb2\ := work.Int.add(\$1646_loop99400_arg\(384 to 415), X"0000000" & X"1");
                    \$1646_loop99400_arg\ := \$1646_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1646_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1646_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1646_loop99400_arg\(32 to 63),32),16), \$1646_loop99400_arg\(64 to 95)) & \$1657_nb2\;
                    state_var607 := \$1646_LOOP99400\;
                  else
                    \$1657_nb2\ := \$1646_loop99400_arg\(384 to 415);
                    \$1646_loop99400_arg\ := \$1646_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1646_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1646_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1646_loop99400_arg\(32 to 63),32),16), \$1646_loop99400_arg\(64 to 95)) & \$1657_nb2\;
                    state_var607 := \$1646_LOOP99400\;
                  end if;
                else
                  \$1646_loop99400_arg\ := \$1646_loop99400_arg\(0 to 31) & \$1646_loop99400_arg\(32 to 63) & 
                  work.Int.add(\$1646_loop99400_arg\(64 to 95), X"0000000" & X"1") & \$1646_loop99400_arg\(96 to 127) & \$1646_loop99400_arg\(128 to 383) & \$1646_loop99400_arg\(384 to 415);
                  state_var607 := \$1646_LOOP99400\;
                end if;
              else
                \$v436\ := work.Int.ge(\$1646_loop99400_arg\(32 to 63), \$1646_loop99400_arg\(0 to 31));
                if \$v436\(0) = '1' then
                  \$1646_loop99400_arg\ := \$1646_loop99400_arg\(0 to 31) & 
                  work.Int.sub(\$1646_loop99400_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1646_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1646_loop99400_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1646_loop99400_arg\(96 to 127) & \$1646_loop99400_arg\(128 to 383) & \$1646_loop99400_arg\(384 to 415);
                  state_var607 := \$1646_LOOP99400\;
                else
                  \$1646_loop99400_result\ := \$1646_loop99400_arg\(384 to 415);
                  \$1607_loop99401_result\ := \$1646_loop99400_result\;
                  \$1599_n\ := \$1607_loop99401_result\;
                  \$1600\ := work.Print.print_string(clk,of_string("rang "));
                  \$1601\ := work.Int.print(clk,\$1598\(1 to 32));
                  \$1602\ := work.Print.print_string(clk,of_string(": "));
                  \$1603\ := work.Int.print(clk,\$1599_n\);
                  \$1606\ := work.Print.print_newline(clk,eclat_unit);
                  \$1604\ := \$1599_n\;
                  \$v423\ := \$$1216_dst_lock\;
                  if \$v423\(0) = '1' then
                    state_var607 := Q_WAIT422;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1597_i\));
                    \$$1216_dst_write\ <= \$1604\; \$$1216_dst_write_request\ <= '1';
                    state_var607 := PAUSE_SET421;
                  end if;
                end if;
              end if;
            when PAR454 =>
              case state_var609 is
              when PAUSE_SET445 =>
                \$$1217_r_write_request\ <= '0';
                release(\$$1217_r_lock\);
                result442 := eclat_unit;
                rdy443 := eclat_true;
                state_var609 := IDLE444;
              when Q_WAIT446 =>
                \$v447\ := \$$1217_r_lock\;
                if \$v447\(0) = '1' then
                  state_var609 := Q_WAIT446;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1597_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var609 := PAUSE_SET445;
                end if;
              when IDLE444 =>
                
              end case;
              
              case state_var608 is
              when PAUSE_GET451 =>
                result448 := \$$1209_src_value\;
                release(\$$1209_src_lock\);
                rdy449 := eclat_true;
                state_var608 := IDLE450;
              when Q_WAIT452 =>
                \$v453\ := \$$1209_src_lock\;
                if \$v453\(0) = '1' then
                  state_var608 := Q_WAIT452;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1597_i\));
                  state_var608 := PAUSE_GET451;
                end if;
              when IDLE450 =>
                
              end case;
              
              \$v455\ := work.Bool.land(rdy443, rdy449);
              if \$v455\(0) = '1' then
                \$1598\ := result442 & result448;
                \$1607_loop99401_id\ := "000000000101";
                \$1607_loop99401_arg\ := X"0000000" & X"2" & X"0000000" & X"1" & X"0000000" & X"1" & eclat_resize(
                work.Vect.infos(256, 48, work.Vect.copy_with(304, 256, 
                                         eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1598\(1 to 32)))(0 to 15),32) & 
                work.Vect.copy_with(304, 256, eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1598\(1 to 32)) & X"0000000" & X"0";
                state_var607 := \$1607_LOOP99401\;
              else
                state_var607 := PAR454;
              end if;
            when PAUSE_GET457 =>
              \$1597_i\ := \$$1217_r_value\;
              release(\$$1217_r_lock\);
              \$v456\ := work.Int.lt(\$1597_i\, std_logic_vector(to_unsigned(\$1209_src\'length,32)));
              if \$v456\(0) = '1' then
                rdy443 := eclat_false;
                \$v447\ := \$$1217_r_lock\;
                if \$v447\(0) = '1' then
                  state_var609 := Q_WAIT446;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1597_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var609 := PAUSE_SET445;
                end if;
                rdy449 := eclat_false;
                \$v453\ := \$$1209_src_lock\;
                if \$v453\(0) = '1' then
                  state_var608 := Q_WAIT452;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1597_i\));
                  state_var608 := PAUSE_GET451;
                end if;
                state_var607 := PAR454;
              else
                \$1594_result\ := eclat_unit;
                result418 := \$1594_result\;
                rdy419 := eclat_true;
                state_var607 := IDLE420;
              end if;
            when PAUSE_SET421 =>
              \$$1216_dst_write_request\ <= '0';
              release(\$$1216_dst_lock\);
              \$1605\ := eclat_unit;
              \$1594_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var607 := \$1594\;
            when Q_WAIT422 =>
              \$v423\ := \$$1216_dst_lock\;
              if \$v423\(0) = '1' then
                state_var607 := Q_WAIT422;
              else
                acquire(\$$1216_dst_lock\);
                \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1597_i\));
                \$$1216_dst_write\ <= \$1604\; \$$1216_dst_write_request\ <= '1';
                state_var607 := PAUSE_SET421;
              end if;
            when Q_WAIT458 =>
              \$v459\ := \$$1217_r_lock\;
              if \$v459\(0) = '1' then
                state_var607 := Q_WAIT458;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var607 := PAUSE_GET457;
              end if;
            when IDLE420 =>
              
            end case;
            
            case state_var604 is
            when \$1660\ =>
              \$v501\ := \$$1217_r_lock\;
              if \$v501\(0) = '1' then
                state_var604 := Q_WAIT500;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var604 := PAUSE_GET499;
              end if;
            when \$1673_LOOP99401\ =>
              \$v481\ := work.Int.le(\$1673_loop99401_arg\(64 to 95), \$1673_loop99401_arg\(96 to 127));
              if \$v481\(0) = '1' then
                \$1683\ := X"0000000" & X"7" & eclat_true;
                \$1682\ := X"0000000" & X"6" & work.Bool.land(""&\$1683\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1683\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1683\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1683\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1683\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1683\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1683\(0 to 31))) & eclat_false)));
                \$1681\ := X"0000000" & X"5" & work.Bool.land(""&\$1682\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1682\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1682\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1682\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1682\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1682\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1682\(0 to 31))) & eclat_false)));
                \$1680\ := X"0000000" & X"4" & work.Bool.land(""&\$1681\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1681\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1681\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1681\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1681\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1681\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1681\(0 to 31))) & eclat_false)));
                \$1679\ := X"0000000" & X"3" & work.Bool.land(""&\$1680\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1680\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1680\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1680\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1680\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1680\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1680\(0 to 31))) & eclat_false)));
                \$1678\ := X"0000000" & X"2" & work.Bool.land(""&\$1679\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1679\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1679\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1679\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1679\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1679\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1679\(0 to 31))) & eclat_false)));
                \$1677\ := X"0000000" & X"1" & work.Bool.land(""&\$1678\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1678\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1678\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1678\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1678\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1678\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1678\(0 to 31))) & eclat_false)));
                \$1676\ := X"0000000" & X"0" & work.Bool.land(""&\$1677\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1677\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1677\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1677\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1677\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1677\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1673_loop99401_arg\(32 to 63), \$1677\(0 to 31))) & eclat_false)));
                \$v475\ := work.Bool.land(""&\$1676\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1676\(0 to 31), X"0000000" & X"1"), \$1673_loop99401_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1676\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1676\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1676\(0 to 31),16),16)), \$1673_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1673_loop99401_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1676\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1673_loop99401_arg\(32 to 63), \$1676\(0 to 31))) & eclat_false)));
                if \$v475\(0) = '1' then
                  \$v470\ := work.Int.eq(work.Int.add(\$1673_loop99401_arg\(32 to 63), X"0000000" & X"1"), \$1673_loop99401_arg\(96 to 127));
                  if \$v470\(0) = '1' then
                    \$1698\ := work.Print.print_string(clk,of_string("foo"));
                    \$1684_nb2\ := work.Int.add(\$1673_loop99401_arg\(384 to 415), X"0000000" & X"1");
                    \$1685_loop99398_id\ := "000000000111";
                    \$1685_loop99398_arg\ := \$1673_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1673_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1673_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1673_loop99401_arg\(32 to 63),32),16), \$1673_loop99401_arg\(64 to 95)) & \$1684_nb2\;
                    state_var604 := \$1685_LOOP99398\;
                  else
                    \$1684_nb2\ := \$1673_loop99401_arg\(384 to 415);
                    \$1685_loop99398_id\ := "000000000111";
                    \$1685_loop99398_arg\ := \$1673_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1673_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1673_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1673_loop99401_arg\(32 to 63),32),16), \$1673_loop99401_arg\(64 to 95)) & \$1684_nb2\;
                    state_var604 := \$1685_LOOP99398\;
                  end if;
                else
                  \$1699_loop99399_id\ := "000000001000";
                  \$1699_loop99399_arg\ := \$1673_loop99401_arg\(0 to 31) & \$1673_loop99401_arg\(32 to 63) & 
                  work.Int.add(\$1673_loop99401_arg\(64 to 95), X"0000000" & X"1") & \$1673_loop99401_arg\(96 to 127) & \$1673_loop99401_arg\(128 to 383) & \$1673_loop99401_arg\(384 to 415);
                  state_var604 := \$1699_LOOP99399\;
                end if;
              else
                \$v480\ := work.Int.ge(\$1673_loop99401_arg\(32 to 63), \$1673_loop99401_arg\(0 to 31));
                if \$v480\(0) = '1' then
                  \$1712_loop99400_id\ := "000000001001";
                  \$1712_loop99400_arg\ := \$1673_loop99401_arg\(0 to 31) & 
                  work.Int.sub(\$1673_loop99401_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1673_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1673_loop99401_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1673_loop99401_arg\(96 to 127) & \$1673_loop99401_arg\(128 to 383) & \$1673_loop99401_arg\(384 to 415);
                  state_var604 := \$1712_LOOP99400\;
                else
                  \$1673_loop99401_result\ := \$1673_loop99401_arg\(384 to 415);
                  \$1665_n\ := \$1673_loop99401_result\;
                  \$1666\ := work.Print.print_string(clk,of_string("rang "));
                  \$1667\ := work.Int.print(clk,\$1664\(1 to 32));
                  \$1668\ := work.Print.print_string(clk,of_string(": "));
                  \$1669\ := work.Int.print(clk,\$1665_n\);
                  \$1672\ := work.Print.print_newline(clk,eclat_unit);
                  \$1670\ := \$1665_n\;
                  \$v465\ := \$$1216_dst_lock\;
                  if \$v465\(0) = '1' then
                    state_var604 := Q_WAIT464;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1663_i\));
                    \$$1216_dst_write\ <= \$1670\; \$$1216_dst_write_request\ <= '1';
                    state_var604 := PAUSE_SET463;
                  end if;
                end if;
              end if;
            when \$1685_LOOP99398\ =>
              \$v469\ := work.Int.le(\$1685_loop99398_arg\(64 to 95), \$1685_loop99398_arg\(96 to 127));
              if \$v469\(0) = '1' then
                \$1695\ := X"0000000" & X"7" & eclat_true;
                \$1694\ := X"0000000" & X"6" & work.Bool.land(""&\$1695\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1695\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1695\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1695\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1695\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1695\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1695\(0 to 31))) & eclat_false)));
                \$1693\ := X"0000000" & X"5" & work.Bool.land(""&\$1694\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1694\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1694\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1694\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1694\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1694\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1694\(0 to 31))) & eclat_false)));
                \$1692\ := X"0000000" & X"4" & work.Bool.land(""&\$1693\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1693\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1693\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1693\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1693\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1693\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1693\(0 to 31))) & eclat_false)));
                \$1691\ := X"0000000" & X"3" & work.Bool.land(""&\$1692\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1692\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1692\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1692\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1692\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1692\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1692\(0 to 31))) & eclat_false)));
                \$1690\ := X"0000000" & X"2" & work.Bool.land(""&\$1691\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1691\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1691\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1691\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1691\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1691\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1691\(0 to 31))) & eclat_false)));
                \$1689\ := X"0000000" & X"1" & work.Bool.land(""&\$1690\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1690\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1690\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1690\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1690\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1690\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1690\(0 to 31))) & eclat_false)));
                \$1688\ := X"0000000" & X"0" & work.Bool.land(""&\$1689\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1689\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1689\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1689\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1689\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1689\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1685_loop99398_arg\(32 to 63), \$1689\(0 to 31))) & eclat_false)));
                \$v467\ := work.Bool.land(""&\$1688\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1688\(0 to 31), X"0000000" & X"1"), \$1685_loop99398_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1688\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1688\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1688\(0 to 31),16),16)), \$1685_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1685_loop99398_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1688\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1685_loop99398_arg\(32 to 63), \$1688\(0 to 31))) & eclat_false)));
                if \$v467\(0) = '1' then
                  \$v466\ := work.Int.eq(work.Int.add(\$1685_loop99398_arg\(32 to 63), X"0000000" & X"1"), \$1685_loop99398_arg\(96 to 127));
                  if \$v466\(0) = '1' then
                    \$1697\ := work.Print.print_string(clk,of_string("foo"));
                    \$1696_nb2\ := work.Int.add(\$1685_loop99398_arg\(384 to 415), X"0000000" & X"1");
                    \$1685_loop99398_arg\ := \$1685_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1685_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1685_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1685_loop99398_arg\(32 to 63),32),16), \$1685_loop99398_arg\(64 to 95)) & \$1696_nb2\;
                    state_var604 := \$1685_LOOP99398\;
                  else
                    \$1696_nb2\ := \$1685_loop99398_arg\(384 to 415);
                    \$1685_loop99398_arg\ := \$1685_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1685_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1685_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1685_loop99398_arg\(32 to 63),32),16), \$1685_loop99398_arg\(64 to 95)) & \$1696_nb2\;
                    state_var604 := \$1685_LOOP99398\;
                  end if;
                else
                  \$1685_loop99398_arg\ := \$1685_loop99398_arg\(0 to 31) & \$1685_loop99398_arg\(32 to 63) & 
                  work.Int.add(\$1685_loop99398_arg\(64 to 95), X"0000000" & X"1") & \$1685_loop99398_arg\(96 to 127) & \$1685_loop99398_arg\(128 to 383) & \$1685_loop99398_arg\(384 to 415);
                  state_var604 := \$1685_LOOP99398\;
                end if;
              else
                \$v468\ := work.Int.ge(\$1685_loop99398_arg\(32 to 63), \$1685_loop99398_arg\(0 to 31));
                if \$v468\(0) = '1' then
                  \$1685_loop99398_arg\ := \$1685_loop99398_arg\(0 to 31) & 
                  work.Int.sub(\$1685_loop99398_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1685_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1685_loop99398_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1685_loop99398_arg\(96 to 127) & \$1685_loop99398_arg\(128 to 383) & \$1685_loop99398_arg\(384 to 415);
                  state_var604 := \$1685_LOOP99398\;
                else
                  \$1685_loop99398_result\ := \$1685_loop99398_arg\(384 to 415);
                  \$1673_loop99401_result\ := \$1685_loop99398_result\;
                  \$1665_n\ := \$1673_loop99401_result\;
                  \$1666\ := work.Print.print_string(clk,of_string("rang "));
                  \$1667\ := work.Int.print(clk,\$1664\(1 to 32));
                  \$1668\ := work.Print.print_string(clk,of_string(": "));
                  \$1669\ := work.Int.print(clk,\$1665_n\);
                  \$1672\ := work.Print.print_newline(clk,eclat_unit);
                  \$1670\ := \$1665_n\;
                  \$v465\ := \$$1216_dst_lock\;
                  if \$v465\(0) = '1' then
                    state_var604 := Q_WAIT464;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1663_i\));
                    \$$1216_dst_write\ <= \$1670\; \$$1216_dst_write_request\ <= '1';
                    state_var604 := PAUSE_SET463;
                  end if;
                end if;
              end if;
            when \$1699_LOOP99399\ =>
              \$v474\ := work.Int.le(\$1699_loop99399_arg\(64 to 95), \$1699_loop99399_arg\(96 to 127));
              if \$v474\(0) = '1' then
                \$1709\ := X"0000000" & X"7" & eclat_true;
                \$1708\ := X"0000000" & X"6" & work.Bool.land(""&\$1709\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1709\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1709\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1709\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1709\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1709\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1709\(0 to 31))) & eclat_false)));
                \$1707\ := X"0000000" & X"5" & work.Bool.land(""&\$1708\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1708\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1708\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1708\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1708\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1708\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1708\(0 to 31))) & eclat_false)));
                \$1706\ := X"0000000" & X"4" & work.Bool.land(""&\$1707\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1707\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1707\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1707\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1707\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1707\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1707\(0 to 31))) & eclat_false)));
                \$1705\ := X"0000000" & X"3" & work.Bool.land(""&\$1706\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1706\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1706\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1706\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1706\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1706\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1706\(0 to 31))) & eclat_false)));
                \$1704\ := X"0000000" & X"2" & work.Bool.land(""&\$1705\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1705\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1705\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1705\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1705\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1705\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1705\(0 to 31))) & eclat_false)));
                \$1703\ := X"0000000" & X"1" & work.Bool.land(""&\$1704\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1704\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1704\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1704\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1704\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1704\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1704\(0 to 31))) & eclat_false)));
                \$1702\ := X"0000000" & X"0" & work.Bool.land(""&\$1703\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1703\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1703\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1703\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1703\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1703\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1699_loop99399_arg\(32 to 63), \$1703\(0 to 31))) & eclat_false)));
                \$v472\ := work.Bool.land(""&\$1702\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1702\(0 to 31), X"0000000" & X"1"), \$1699_loop99399_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1702\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1702\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1702\(0 to 31),16),16)), \$1699_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1699_loop99399_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1702\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1699_loop99399_arg\(32 to 63), \$1702\(0 to 31))) & eclat_false)));
                if \$v472\(0) = '1' then
                  \$v471\ := work.Int.eq(work.Int.add(\$1699_loop99399_arg\(32 to 63), X"0000000" & X"1"), \$1699_loop99399_arg\(96 to 127));
                  if \$v471\(0) = '1' then
                    \$1711\ := work.Print.print_string(clk,of_string("foo"));
                    \$1710_nb2\ := work.Int.add(\$1699_loop99399_arg\(384 to 415), X"0000000" & X"1");
                    \$1699_loop99399_arg\ := \$1699_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1699_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1699_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1699_loop99399_arg\(32 to 63),32),16), \$1699_loop99399_arg\(64 to 95)) & \$1710_nb2\;
                    state_var604 := \$1699_LOOP99399\;
                  else
                    \$1710_nb2\ := \$1699_loop99399_arg\(384 to 415);
                    \$1699_loop99399_arg\ := \$1699_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1699_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1699_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1699_loop99399_arg\(32 to 63),32),16), \$1699_loop99399_arg\(64 to 95)) & \$1710_nb2\;
                    state_var604 := \$1699_LOOP99399\;
                  end if;
                else
                  \$1699_loop99399_arg\ := \$1699_loop99399_arg\(0 to 31) & \$1699_loop99399_arg\(32 to 63) & 
                  work.Int.add(\$1699_loop99399_arg\(64 to 95), X"0000000" & X"1") & \$1699_loop99399_arg\(96 to 127) & \$1699_loop99399_arg\(128 to 383) & \$1699_loop99399_arg\(384 to 415);
                  state_var604 := \$1699_LOOP99399\;
                end if;
              else
                \$v473\ := work.Int.ge(\$1699_loop99399_arg\(32 to 63), \$1699_loop99399_arg\(0 to 31));
                if \$v473\(0) = '1' then
                  \$1699_loop99399_arg\ := \$1699_loop99399_arg\(0 to 31) & 
                  work.Int.sub(\$1699_loop99399_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1699_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1699_loop99399_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1699_loop99399_arg\(96 to 127) & \$1699_loop99399_arg\(128 to 383) & \$1699_loop99399_arg\(384 to 415);
                  state_var604 := \$1699_LOOP99399\;
                else
                  \$1699_loop99399_result\ := \$1699_loop99399_arg\(384 to 415);
                  \$1673_loop99401_result\ := \$1699_loop99399_result\;
                  \$1665_n\ := \$1673_loop99401_result\;
                  \$1666\ := work.Print.print_string(clk,of_string("rang "));
                  \$1667\ := work.Int.print(clk,\$1664\(1 to 32));
                  \$1668\ := work.Print.print_string(clk,of_string(": "));
                  \$1669\ := work.Int.print(clk,\$1665_n\);
                  \$1672\ := work.Print.print_newline(clk,eclat_unit);
                  \$1670\ := \$1665_n\;
                  \$v465\ := \$$1216_dst_lock\;
                  if \$v465\(0) = '1' then
                    state_var604 := Q_WAIT464;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1663_i\));
                    \$$1216_dst_write\ <= \$1670\; \$$1216_dst_write_request\ <= '1';
                    state_var604 := PAUSE_SET463;
                  end if;
                end if;
              end if;
            when \$1712_LOOP99400\ =>
              \$v479\ := work.Int.le(\$1712_loop99400_arg\(64 to 95), \$1712_loop99400_arg\(96 to 127));
              if \$v479\(0) = '1' then
                \$1722\ := X"0000000" & X"7" & eclat_true;
                \$1721\ := X"0000000" & X"6" & work.Bool.land(""&\$1722\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1722\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1722\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1722\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1722\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1722\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1722\(0 to 31))) & eclat_false)));
                \$1720\ := X"0000000" & X"5" & work.Bool.land(""&\$1721\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1721\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1721\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1721\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1721\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1721\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1721\(0 to 31))) & eclat_false)));
                \$1719\ := X"0000000" & X"4" & work.Bool.land(""&\$1720\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1720\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1720\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1720\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1720\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1720\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1720\(0 to 31))) & eclat_false)));
                \$1718\ := X"0000000" & X"3" & work.Bool.land(""&\$1719\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1719\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1719\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1719\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1719\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1719\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1719\(0 to 31))) & eclat_false)));
                \$1717\ := X"0000000" & X"2" & work.Bool.land(""&\$1718\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1718\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1718\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1718\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1718\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1718\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1718\(0 to 31))) & eclat_false)));
                \$1716\ := X"0000000" & X"1" & work.Bool.land(""&\$1717\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1717\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1717\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1717\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1717\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1717\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1717\(0 to 31))) & eclat_false)));
                \$1715\ := X"0000000" & X"0" & work.Bool.land(""&\$1716\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1716\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1716\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1716\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1716\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1716\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1712_loop99400_arg\(32 to 63), \$1716\(0 to 31))) & eclat_false)));
                \$v477\ := work.Bool.land(""&\$1715\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1715\(0 to 31), X"0000000" & X"1"), \$1712_loop99400_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1715\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1715\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1715\(0 to 31),16),16)), \$1712_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1712_loop99400_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1715\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1712_loop99400_arg\(32 to 63), \$1715\(0 to 31))) & eclat_false)));
                if \$v477\(0) = '1' then
                  \$v476\ := work.Int.eq(work.Int.add(\$1712_loop99400_arg\(32 to 63), X"0000000" & X"1"), \$1712_loop99400_arg\(96 to 127));
                  if \$v476\(0) = '1' then
                    \$1724\ := work.Print.print_string(clk,of_string("foo"));
                    \$1723_nb2\ := work.Int.add(\$1712_loop99400_arg\(384 to 415), X"0000000" & X"1");
                    \$1712_loop99400_arg\ := \$1712_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1712_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1712_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1712_loop99400_arg\(32 to 63),32),16), \$1712_loop99400_arg\(64 to 95)) & \$1723_nb2\;
                    state_var604 := \$1712_LOOP99400\;
                  else
                    \$1723_nb2\ := \$1712_loop99400_arg\(384 to 415);
                    \$1712_loop99400_arg\ := \$1712_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1712_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1712_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1712_loop99400_arg\(32 to 63),32),16), \$1712_loop99400_arg\(64 to 95)) & \$1723_nb2\;
                    state_var604 := \$1712_LOOP99400\;
                  end if;
                else
                  \$1712_loop99400_arg\ := \$1712_loop99400_arg\(0 to 31) & \$1712_loop99400_arg\(32 to 63) & 
                  work.Int.add(\$1712_loop99400_arg\(64 to 95), X"0000000" & X"1") & \$1712_loop99400_arg\(96 to 127) & \$1712_loop99400_arg\(128 to 383) & \$1712_loop99400_arg\(384 to 415);
                  state_var604 := \$1712_LOOP99400\;
                end if;
              else
                \$v478\ := work.Int.ge(\$1712_loop99400_arg\(32 to 63), \$1712_loop99400_arg\(0 to 31));
                if \$v478\(0) = '1' then
                  \$1712_loop99400_arg\ := \$1712_loop99400_arg\(0 to 31) & 
                  work.Int.sub(\$1712_loop99400_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1712_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1712_loop99400_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1712_loop99400_arg\(96 to 127) & \$1712_loop99400_arg\(128 to 383) & \$1712_loop99400_arg\(384 to 415);
                  state_var604 := \$1712_LOOP99400\;
                else
                  \$1712_loop99400_result\ := \$1712_loop99400_arg\(384 to 415);
                  \$1673_loop99401_result\ := \$1712_loop99400_result\;
                  \$1665_n\ := \$1673_loop99401_result\;
                  \$1666\ := work.Print.print_string(clk,of_string("rang "));
                  \$1667\ := work.Int.print(clk,\$1664\(1 to 32));
                  \$1668\ := work.Print.print_string(clk,of_string(": "));
                  \$1669\ := work.Int.print(clk,\$1665_n\);
                  \$1672\ := work.Print.print_newline(clk,eclat_unit);
                  \$1670\ := \$1665_n\;
                  \$v465\ := \$$1216_dst_lock\;
                  if \$v465\(0) = '1' then
                    state_var604 := Q_WAIT464;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1663_i\));
                    \$$1216_dst_write\ <= \$1670\; \$$1216_dst_write_request\ <= '1';
                    state_var604 := PAUSE_SET463;
                  end if;
                end if;
              end if;
            when PAR496 =>
              case state_var606 is
              when PAUSE_SET487 =>
                \$$1217_r_write_request\ <= '0';
                release(\$$1217_r_lock\);
                result484 := eclat_unit;
                rdy485 := eclat_true;
                state_var606 := IDLE486;
              when Q_WAIT488 =>
                \$v489\ := \$$1217_r_lock\;
                if \$v489\(0) = '1' then
                  state_var606 := Q_WAIT488;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1663_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var606 := PAUSE_SET487;
                end if;
              when IDLE486 =>
                
              end case;
              
              case state_var605 is
              when PAUSE_GET493 =>
                result490 := \$$1209_src_value\;
                release(\$$1209_src_lock\);
                rdy491 := eclat_true;
                state_var605 := IDLE492;
              when Q_WAIT494 =>
                \$v495\ := \$$1209_src_lock\;
                if \$v495\(0) = '1' then
                  state_var605 := Q_WAIT494;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1663_i\));
                  state_var605 := PAUSE_GET493;
                end if;
              when IDLE492 =>
                
              end case;
              
              \$v497\ := work.Bool.land(rdy485, rdy491);
              if \$v497\(0) = '1' then
                \$1664\ := result484 & result490;
                \$1673_loop99401_id\ := "000000001010";
                \$1673_loop99401_arg\ := X"0000000" & X"2" & X"0000000" & X"1" & X"0000000" & X"1" & eclat_resize(
                work.Vect.infos(256, 48, work.Vect.copy_with(304, 256, 
                                         eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1664\(1 to 32)))(0 to 15),32) & 
                work.Vect.copy_with(304, 256, eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1664\(1 to 32)) & X"0000000" & X"0";
                state_var604 := \$1673_LOOP99401\;
              else
                state_var604 := PAR496;
              end if;
            when PAUSE_GET499 =>
              \$1663_i\ := \$$1217_r_value\;
              release(\$$1217_r_lock\);
              \$v498\ := work.Int.lt(\$1663_i\, std_logic_vector(to_unsigned(\$1209_src\'length,32)));
              if \$v498\(0) = '1' then
                rdy485 := eclat_false;
                \$v489\ := \$$1217_r_lock\;
                if \$v489\(0) = '1' then
                  state_var606 := Q_WAIT488;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1663_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var606 := PAUSE_SET487;
                end if;
                rdy491 := eclat_false;
                \$v495\ := \$$1209_src_lock\;
                if \$v495\(0) = '1' then
                  state_var605 := Q_WAIT494;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1663_i\));
                  state_var605 := PAUSE_GET493;
                end if;
                state_var604 := PAR496;
              else
                \$1660_result\ := eclat_unit;
                result460 := \$1660_result\;
                rdy461 := eclat_true;
                state_var604 := IDLE462;
              end if;
            when PAUSE_SET463 =>
              \$$1216_dst_write_request\ <= '0';
              release(\$$1216_dst_lock\);
              \$1671\ := eclat_unit;
              \$1660_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var604 := \$1660\;
            when Q_WAIT464 =>
              \$v465\ := \$$1216_dst_lock\;
              if \$v465\(0) = '1' then
                state_var604 := Q_WAIT464;
              else
                acquire(\$$1216_dst_lock\);
                \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1663_i\));
                \$$1216_dst_write\ <= \$1670\; \$$1216_dst_write_request\ <= '1';
                state_var604 := PAUSE_SET463;
              end if;
            when Q_WAIT500 =>
              \$v501\ := \$$1217_r_lock\;
              if \$v501\(0) = '1' then
                state_var604 := Q_WAIT500;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var604 := PAUSE_GET499;
              end if;
            when IDLE462 =>
              
            end case;
            
            case state_var601 is
            when \$1726\ =>
              \$v543\ := \$$1217_r_lock\;
              if \$v543\(0) = '1' then
                state_var601 := Q_WAIT542;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var601 := PAUSE_GET541;
              end if;
            when \$1739_LOOP99401\ =>
              \$v523\ := work.Int.le(\$1739_loop99401_arg\(64 to 95), \$1739_loop99401_arg\(96 to 127));
              if \$v523\(0) = '1' then
                \$1749\ := X"0000000" & X"7" & eclat_true;
                \$1748\ := X"0000000" & X"6" & work.Bool.land(""&\$1749\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1749\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1749\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1749\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1749\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1749\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1749\(0 to 31))) & eclat_false)));
                \$1747\ := X"0000000" & X"5" & work.Bool.land(""&\$1748\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1748\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1748\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1748\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1748\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1748\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1748\(0 to 31))) & eclat_false)));
                \$1746\ := X"0000000" & X"4" & work.Bool.land(""&\$1747\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1747\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1747\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1747\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1747\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1747\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1747\(0 to 31))) & eclat_false)));
                \$1745\ := X"0000000" & X"3" & work.Bool.land(""&\$1746\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1746\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1746\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1746\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1746\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1746\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1746\(0 to 31))) & eclat_false)));
                \$1744\ := X"0000000" & X"2" & work.Bool.land(""&\$1745\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1745\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1745\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1745\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1745\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1745\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1745\(0 to 31))) & eclat_false)));
                \$1743\ := X"0000000" & X"1" & work.Bool.land(""&\$1744\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1744\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1744\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1744\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1744\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1744\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1744\(0 to 31))) & eclat_false)));
                \$1742\ := X"0000000" & X"0" & work.Bool.land(""&\$1743\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1743\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1743\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1743\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1743\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1743\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1739_loop99401_arg\(32 to 63), \$1743\(0 to 31))) & eclat_false)));
                \$v517\ := work.Bool.land(""&\$1742\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1742\(0 to 31), X"0000000" & X"1"), \$1739_loop99401_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1742\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1742\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1742\(0 to 31),16),16)), \$1739_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1739_loop99401_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1742\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1739_loop99401_arg\(32 to 63), \$1742\(0 to 31))) & eclat_false)));
                if \$v517\(0) = '1' then
                  \$v512\ := work.Int.eq(work.Int.add(\$1739_loop99401_arg\(32 to 63), X"0000000" & X"1"), \$1739_loop99401_arg\(96 to 127));
                  if \$v512\(0) = '1' then
                    \$1764\ := work.Print.print_string(clk,of_string("foo"));
                    \$1750_nb2\ := work.Int.add(\$1739_loop99401_arg\(384 to 415), X"0000000" & X"1");
                    \$1751_loop99398_id\ := "000000001100";
                    \$1751_loop99398_arg\ := \$1739_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1739_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1739_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1739_loop99401_arg\(32 to 63),32),16), \$1739_loop99401_arg\(64 to 95)) & \$1750_nb2\;
                    state_var601 := \$1751_LOOP99398\;
                  else
                    \$1750_nb2\ := \$1739_loop99401_arg\(384 to 415);
                    \$1751_loop99398_id\ := "000000001100";
                    \$1751_loop99398_arg\ := \$1739_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1739_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1739_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1739_loop99401_arg\(32 to 63),32),16), \$1739_loop99401_arg\(64 to 95)) & \$1750_nb2\;
                    state_var601 := \$1751_LOOP99398\;
                  end if;
                else
                  \$1765_loop99399_id\ := "000000001101";
                  \$1765_loop99399_arg\ := \$1739_loop99401_arg\(0 to 31) & \$1739_loop99401_arg\(32 to 63) & 
                  work.Int.add(\$1739_loop99401_arg\(64 to 95), X"0000000" & X"1") & \$1739_loop99401_arg\(96 to 127) & \$1739_loop99401_arg\(128 to 383) & \$1739_loop99401_arg\(384 to 415);
                  state_var601 := \$1765_LOOP99399\;
                end if;
              else
                \$v522\ := work.Int.ge(\$1739_loop99401_arg\(32 to 63), \$1739_loop99401_arg\(0 to 31));
                if \$v522\(0) = '1' then
                  \$1778_loop99400_id\ := "000000001110";
                  \$1778_loop99400_arg\ := \$1739_loop99401_arg\(0 to 31) & 
                  work.Int.sub(\$1739_loop99401_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1739_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1739_loop99401_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1739_loop99401_arg\(96 to 127) & \$1739_loop99401_arg\(128 to 383) & \$1739_loop99401_arg\(384 to 415);
                  state_var601 := \$1778_LOOP99400\;
                else
                  \$1739_loop99401_result\ := \$1739_loop99401_arg\(384 to 415);
                  \$1731_n\ := \$1739_loop99401_result\;
                  \$1732\ := work.Print.print_string(clk,of_string("rang "));
                  \$1733\ := work.Int.print(clk,\$1730\(1 to 32));
                  \$1734\ := work.Print.print_string(clk,of_string(": "));
                  \$1735\ := work.Int.print(clk,\$1731_n\);
                  \$1738\ := work.Print.print_newline(clk,eclat_unit);
                  \$1736\ := \$1731_n\;
                  \$v507\ := \$$1216_dst_lock\;
                  if \$v507\(0) = '1' then
                    state_var601 := Q_WAIT506;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1729_i\));
                    \$$1216_dst_write\ <= \$1736\; \$$1216_dst_write_request\ <= '1';
                    state_var601 := PAUSE_SET505;
                  end if;
                end if;
              end if;
            when \$1751_LOOP99398\ =>
              \$v511\ := work.Int.le(\$1751_loop99398_arg\(64 to 95), \$1751_loop99398_arg\(96 to 127));
              if \$v511\(0) = '1' then
                \$1761\ := X"0000000" & X"7" & eclat_true;
                \$1760\ := X"0000000" & X"6" & work.Bool.land(""&\$1761\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1761\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1761\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1761\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1761\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1761\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1761\(0 to 31))) & eclat_false)));
                \$1759\ := X"0000000" & X"5" & work.Bool.land(""&\$1760\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1760\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1760\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1760\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1760\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1760\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1760\(0 to 31))) & eclat_false)));
                \$1758\ := X"0000000" & X"4" & work.Bool.land(""&\$1759\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1759\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1759\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1759\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1759\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1759\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1759\(0 to 31))) & eclat_false)));
                \$1757\ := X"0000000" & X"3" & work.Bool.land(""&\$1758\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1758\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1758\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1758\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1758\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1758\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1758\(0 to 31))) & eclat_false)));
                \$1756\ := X"0000000" & X"2" & work.Bool.land(""&\$1757\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1757\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1757\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1757\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1757\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1757\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1757\(0 to 31))) & eclat_false)));
                \$1755\ := X"0000000" & X"1" & work.Bool.land(""&\$1756\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1756\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1756\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1756\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1756\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1756\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1756\(0 to 31))) & eclat_false)));
                \$1754\ := X"0000000" & X"0" & work.Bool.land(""&\$1755\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1755\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1755\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1755\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1755\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1755\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1751_loop99398_arg\(32 to 63), \$1755\(0 to 31))) & eclat_false)));
                \$v509\ := work.Bool.land(""&\$1754\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1754\(0 to 31), X"0000000" & X"1"), \$1751_loop99398_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1754\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1754\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1754\(0 to 31),16),16)), \$1751_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1751_loop99398_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1754\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1751_loop99398_arg\(32 to 63), \$1754\(0 to 31))) & eclat_false)));
                if \$v509\(0) = '1' then
                  \$v508\ := work.Int.eq(work.Int.add(\$1751_loop99398_arg\(32 to 63), X"0000000" & X"1"), \$1751_loop99398_arg\(96 to 127));
                  if \$v508\(0) = '1' then
                    \$1763\ := work.Print.print_string(clk,of_string("foo"));
                    \$1762_nb2\ := work.Int.add(\$1751_loop99398_arg\(384 to 415), X"0000000" & X"1");
                    \$1751_loop99398_arg\ := \$1751_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1751_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1751_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1751_loop99398_arg\(32 to 63),32),16), \$1751_loop99398_arg\(64 to 95)) & \$1762_nb2\;
                    state_var601 := \$1751_LOOP99398\;
                  else
                    \$1762_nb2\ := \$1751_loop99398_arg\(384 to 415);
                    \$1751_loop99398_arg\ := \$1751_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1751_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1751_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1751_loop99398_arg\(32 to 63),32),16), \$1751_loop99398_arg\(64 to 95)) & \$1762_nb2\;
                    state_var601 := \$1751_LOOP99398\;
                  end if;
                else
                  \$1751_loop99398_arg\ := \$1751_loop99398_arg\(0 to 31) & \$1751_loop99398_arg\(32 to 63) & 
                  work.Int.add(\$1751_loop99398_arg\(64 to 95), X"0000000" & X"1") & \$1751_loop99398_arg\(96 to 127) & \$1751_loop99398_arg\(128 to 383) & \$1751_loop99398_arg\(384 to 415);
                  state_var601 := \$1751_LOOP99398\;
                end if;
              else
                \$v510\ := work.Int.ge(\$1751_loop99398_arg\(32 to 63), \$1751_loop99398_arg\(0 to 31));
                if \$v510\(0) = '1' then
                  \$1751_loop99398_arg\ := \$1751_loop99398_arg\(0 to 31) & 
                  work.Int.sub(\$1751_loop99398_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1751_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1751_loop99398_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1751_loop99398_arg\(96 to 127) & \$1751_loop99398_arg\(128 to 383) & \$1751_loop99398_arg\(384 to 415);
                  state_var601 := \$1751_LOOP99398\;
                else
                  \$1751_loop99398_result\ := \$1751_loop99398_arg\(384 to 415);
                  \$1739_loop99401_result\ := \$1751_loop99398_result\;
                  \$1731_n\ := \$1739_loop99401_result\;
                  \$1732\ := work.Print.print_string(clk,of_string("rang "));
                  \$1733\ := work.Int.print(clk,\$1730\(1 to 32));
                  \$1734\ := work.Print.print_string(clk,of_string(": "));
                  \$1735\ := work.Int.print(clk,\$1731_n\);
                  \$1738\ := work.Print.print_newline(clk,eclat_unit);
                  \$1736\ := \$1731_n\;
                  \$v507\ := \$$1216_dst_lock\;
                  if \$v507\(0) = '1' then
                    state_var601 := Q_WAIT506;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1729_i\));
                    \$$1216_dst_write\ <= \$1736\; \$$1216_dst_write_request\ <= '1';
                    state_var601 := PAUSE_SET505;
                  end if;
                end if;
              end if;
            when \$1765_LOOP99399\ =>
              \$v516\ := work.Int.le(\$1765_loop99399_arg\(64 to 95), \$1765_loop99399_arg\(96 to 127));
              if \$v516\(0) = '1' then
                \$1775\ := X"0000000" & X"7" & eclat_true;
                \$1774\ := X"0000000" & X"6" & work.Bool.land(""&\$1775\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1775\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1775\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1775\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1775\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1775\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1775\(0 to 31))) & eclat_false)));
                \$1773\ := X"0000000" & X"5" & work.Bool.land(""&\$1774\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1774\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1774\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1774\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1774\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1774\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1774\(0 to 31))) & eclat_false)));
                \$1772\ := X"0000000" & X"4" & work.Bool.land(""&\$1773\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1773\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1773\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1773\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1773\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1773\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1773\(0 to 31))) & eclat_false)));
                \$1771\ := X"0000000" & X"3" & work.Bool.land(""&\$1772\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1772\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1772\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1772\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1772\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1772\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1772\(0 to 31))) & eclat_false)));
                \$1770\ := X"0000000" & X"2" & work.Bool.land(""&\$1771\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1771\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1771\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1771\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1771\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1771\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1771\(0 to 31))) & eclat_false)));
                \$1769\ := X"0000000" & X"1" & work.Bool.land(""&\$1770\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1770\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1770\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1770\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1770\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1770\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1770\(0 to 31))) & eclat_false)));
                \$1768\ := X"0000000" & X"0" & work.Bool.land(""&\$1769\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1769\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1769\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1769\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1769\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1769\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1765_loop99399_arg\(32 to 63), \$1769\(0 to 31))) & eclat_false)));
                \$v514\ := work.Bool.land(""&\$1768\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1768\(0 to 31), X"0000000" & X"1"), \$1765_loop99399_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1768\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1768\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1768\(0 to 31),16),16)), \$1765_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1765_loop99399_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1768\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1765_loop99399_arg\(32 to 63), \$1768\(0 to 31))) & eclat_false)));
                if \$v514\(0) = '1' then
                  \$v513\ := work.Int.eq(work.Int.add(\$1765_loop99399_arg\(32 to 63), X"0000000" & X"1"), \$1765_loop99399_arg\(96 to 127));
                  if \$v513\(0) = '1' then
                    \$1777\ := work.Print.print_string(clk,of_string("foo"));
                    \$1776_nb2\ := work.Int.add(\$1765_loop99399_arg\(384 to 415), X"0000000" & X"1");
                    \$1765_loop99399_arg\ := \$1765_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1765_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1765_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1765_loop99399_arg\(32 to 63),32),16), \$1765_loop99399_arg\(64 to 95)) & \$1776_nb2\;
                    state_var601 := \$1765_LOOP99399\;
                  else
                    \$1776_nb2\ := \$1765_loop99399_arg\(384 to 415);
                    \$1765_loop99399_arg\ := \$1765_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1765_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1765_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1765_loop99399_arg\(32 to 63),32),16), \$1765_loop99399_arg\(64 to 95)) & \$1776_nb2\;
                    state_var601 := \$1765_LOOP99399\;
                  end if;
                else
                  \$1765_loop99399_arg\ := \$1765_loop99399_arg\(0 to 31) & \$1765_loop99399_arg\(32 to 63) & 
                  work.Int.add(\$1765_loop99399_arg\(64 to 95), X"0000000" & X"1") & \$1765_loop99399_arg\(96 to 127) & \$1765_loop99399_arg\(128 to 383) & \$1765_loop99399_arg\(384 to 415);
                  state_var601 := \$1765_LOOP99399\;
                end if;
              else
                \$v515\ := work.Int.ge(\$1765_loop99399_arg\(32 to 63), \$1765_loop99399_arg\(0 to 31));
                if \$v515\(0) = '1' then
                  \$1765_loop99399_arg\ := \$1765_loop99399_arg\(0 to 31) & 
                  work.Int.sub(\$1765_loop99399_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1765_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1765_loop99399_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1765_loop99399_arg\(96 to 127) & \$1765_loop99399_arg\(128 to 383) & \$1765_loop99399_arg\(384 to 415);
                  state_var601 := \$1765_LOOP99399\;
                else
                  \$1765_loop99399_result\ := \$1765_loop99399_arg\(384 to 415);
                  \$1739_loop99401_result\ := \$1765_loop99399_result\;
                  \$1731_n\ := \$1739_loop99401_result\;
                  \$1732\ := work.Print.print_string(clk,of_string("rang "));
                  \$1733\ := work.Int.print(clk,\$1730\(1 to 32));
                  \$1734\ := work.Print.print_string(clk,of_string(": "));
                  \$1735\ := work.Int.print(clk,\$1731_n\);
                  \$1738\ := work.Print.print_newline(clk,eclat_unit);
                  \$1736\ := \$1731_n\;
                  \$v507\ := \$$1216_dst_lock\;
                  if \$v507\(0) = '1' then
                    state_var601 := Q_WAIT506;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1729_i\));
                    \$$1216_dst_write\ <= \$1736\; \$$1216_dst_write_request\ <= '1';
                    state_var601 := PAUSE_SET505;
                  end if;
                end if;
              end if;
            when \$1778_LOOP99400\ =>
              \$v521\ := work.Int.le(\$1778_loop99400_arg\(64 to 95), \$1778_loop99400_arg\(96 to 127));
              if \$v521\(0) = '1' then
                \$1788\ := X"0000000" & X"7" & eclat_true;
                \$1787\ := X"0000000" & X"6" & work.Bool.land(""&\$1788\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1788\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1788\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1788\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1788\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1788\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1788\(0 to 31))) & eclat_false)));
                \$1786\ := X"0000000" & X"5" & work.Bool.land(""&\$1787\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1787\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1787\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1787\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1787\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1787\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1787\(0 to 31))) & eclat_false)));
                \$1785\ := X"0000000" & X"4" & work.Bool.land(""&\$1786\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1786\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1786\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1786\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1786\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1786\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1786\(0 to 31))) & eclat_false)));
                \$1784\ := X"0000000" & X"3" & work.Bool.land(""&\$1785\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1785\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1785\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1785\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1785\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1785\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1785\(0 to 31))) & eclat_false)));
                \$1783\ := X"0000000" & X"2" & work.Bool.land(""&\$1784\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1784\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1784\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1784\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1784\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1784\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1784\(0 to 31))) & eclat_false)));
                \$1782\ := X"0000000" & X"1" & work.Bool.land(""&\$1783\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1783\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1783\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1783\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1783\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1783\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1783\(0 to 31))) & eclat_false)));
                \$1781\ := X"0000000" & X"0" & work.Bool.land(""&\$1782\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1782\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1782\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1782\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1782\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1782\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1778_loop99400_arg\(32 to 63), \$1782\(0 to 31))) & eclat_false)));
                \$v519\ := work.Bool.land(""&\$1781\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1781\(0 to 31), X"0000000" & X"1"), \$1778_loop99400_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1781\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1781\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1781\(0 to 31),16),16)), \$1778_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1778_loop99400_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1781\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1778_loop99400_arg\(32 to 63), \$1781\(0 to 31))) & eclat_false)));
                if \$v519\(0) = '1' then
                  \$v518\ := work.Int.eq(work.Int.add(\$1778_loop99400_arg\(32 to 63), X"0000000" & X"1"), \$1778_loop99400_arg\(96 to 127));
                  if \$v518\(0) = '1' then
                    \$1790\ := work.Print.print_string(clk,of_string("foo"));
                    \$1789_nb2\ := work.Int.add(\$1778_loop99400_arg\(384 to 415), X"0000000" & X"1");
                    \$1778_loop99400_arg\ := \$1778_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1778_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1778_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1778_loop99400_arg\(32 to 63),32),16), \$1778_loop99400_arg\(64 to 95)) & \$1789_nb2\;
                    state_var601 := \$1778_LOOP99400\;
                  else
                    \$1789_nb2\ := \$1778_loop99400_arg\(384 to 415);
                    \$1778_loop99400_arg\ := \$1778_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1778_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1778_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1778_loop99400_arg\(32 to 63),32),16), \$1778_loop99400_arg\(64 to 95)) & \$1789_nb2\;
                    state_var601 := \$1778_LOOP99400\;
                  end if;
                else
                  \$1778_loop99400_arg\ := \$1778_loop99400_arg\(0 to 31) & \$1778_loop99400_arg\(32 to 63) & 
                  work.Int.add(\$1778_loop99400_arg\(64 to 95), X"0000000" & X"1") & \$1778_loop99400_arg\(96 to 127) & \$1778_loop99400_arg\(128 to 383) & \$1778_loop99400_arg\(384 to 415);
                  state_var601 := \$1778_LOOP99400\;
                end if;
              else
                \$v520\ := work.Int.ge(\$1778_loop99400_arg\(32 to 63), \$1778_loop99400_arg\(0 to 31));
                if \$v520\(0) = '1' then
                  \$1778_loop99400_arg\ := \$1778_loop99400_arg\(0 to 31) & 
                  work.Int.sub(\$1778_loop99400_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1778_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1778_loop99400_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1778_loop99400_arg\(96 to 127) & \$1778_loop99400_arg\(128 to 383) & \$1778_loop99400_arg\(384 to 415);
                  state_var601 := \$1778_LOOP99400\;
                else
                  \$1778_loop99400_result\ := \$1778_loop99400_arg\(384 to 415);
                  \$1739_loop99401_result\ := \$1778_loop99400_result\;
                  \$1731_n\ := \$1739_loop99401_result\;
                  \$1732\ := work.Print.print_string(clk,of_string("rang "));
                  \$1733\ := work.Int.print(clk,\$1730\(1 to 32));
                  \$1734\ := work.Print.print_string(clk,of_string(": "));
                  \$1735\ := work.Int.print(clk,\$1731_n\);
                  \$1738\ := work.Print.print_newline(clk,eclat_unit);
                  \$1736\ := \$1731_n\;
                  \$v507\ := \$$1216_dst_lock\;
                  if \$v507\(0) = '1' then
                    state_var601 := Q_WAIT506;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1729_i\));
                    \$$1216_dst_write\ <= \$1736\; \$$1216_dst_write_request\ <= '1';
                    state_var601 := PAUSE_SET505;
                  end if;
                end if;
              end if;
            when PAR538 =>
              case state_var603 is
              when PAUSE_SET529 =>
                \$$1217_r_write_request\ <= '0';
                release(\$$1217_r_lock\);
                result526 := eclat_unit;
                rdy527 := eclat_true;
                state_var603 := IDLE528;
              when Q_WAIT530 =>
                \$v531\ := \$$1217_r_lock\;
                if \$v531\(0) = '1' then
                  state_var603 := Q_WAIT530;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1729_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var603 := PAUSE_SET529;
                end if;
              when IDLE528 =>
                
              end case;
              
              case state_var602 is
              when PAUSE_GET535 =>
                result532 := \$$1209_src_value\;
                release(\$$1209_src_lock\);
                rdy533 := eclat_true;
                state_var602 := IDLE534;
              when Q_WAIT536 =>
                \$v537\ := \$$1209_src_lock\;
                if \$v537\(0) = '1' then
                  state_var602 := Q_WAIT536;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1729_i\));
                  state_var602 := PAUSE_GET535;
                end if;
              when IDLE534 =>
                
              end case;
              
              \$v539\ := work.Bool.land(rdy527, rdy533);
              if \$v539\(0) = '1' then
                \$1730\ := result526 & result532;
                \$1739_loop99401_id\ := "000000001111";
                \$1739_loop99401_arg\ := X"0000000" & X"2" & X"0000000" & X"1" & X"0000000" & X"1" & eclat_resize(
                work.Vect.infos(256, 48, work.Vect.copy_with(304, 256, 
                                         eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1730\(1 to 32)))(0 to 15),32) & 
                work.Vect.copy_with(304, 256, eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1730\(1 to 32)) & X"0000000" & X"0";
                state_var601 := \$1739_LOOP99401\;
              else
                state_var601 := PAR538;
              end if;
            when PAUSE_GET541 =>
              \$1729_i\ := \$$1217_r_value\;
              release(\$$1217_r_lock\);
              \$v540\ := work.Int.lt(\$1729_i\, std_logic_vector(to_unsigned(\$1209_src\'length,32)));
              if \$v540\(0) = '1' then
                rdy527 := eclat_false;
                \$v531\ := \$$1217_r_lock\;
                if \$v531\(0) = '1' then
                  state_var603 := Q_WAIT530;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1729_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var603 := PAUSE_SET529;
                end if;
                rdy533 := eclat_false;
                \$v537\ := \$$1209_src_lock\;
                if \$v537\(0) = '1' then
                  state_var602 := Q_WAIT536;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1729_i\));
                  state_var602 := PAUSE_GET535;
                end if;
                state_var601 := PAR538;
              else
                \$1726_result\ := eclat_unit;
                result502 := \$1726_result\;
                rdy503 := eclat_true;
                state_var601 := IDLE504;
              end if;
            when PAUSE_SET505 =>
              \$$1216_dst_write_request\ <= '0';
              release(\$$1216_dst_lock\);
              \$1737\ := eclat_unit;
              \$1726_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var601 := \$1726\;
            when Q_WAIT506 =>
              \$v507\ := \$$1216_dst_lock\;
              if \$v507\(0) = '1' then
                state_var601 := Q_WAIT506;
              else
                acquire(\$$1216_dst_lock\);
                \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1729_i\));
                \$$1216_dst_write\ <= \$1736\; \$$1216_dst_write_request\ <= '1';
                state_var601 := PAUSE_SET505;
              end if;
            when Q_WAIT542 =>
              \$v543\ := \$$1217_r_lock\;
              if \$v543\(0) = '1' then
                state_var601 := Q_WAIT542;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var601 := PAUSE_GET541;
              end if;
            when IDLE504 =>
              
            end case;
            
            case state_var598 is
            when \$1792\ =>
              \$v585\ := \$$1217_r_lock\;
              if \$v585\(0) = '1' then
                state_var598 := Q_WAIT584;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var598 := PAUSE_GET583;
              end if;
            when \$1805_LOOP99401\ =>
              \$v565\ := work.Int.le(\$1805_loop99401_arg\(64 to 95), \$1805_loop99401_arg\(96 to 127));
              if \$v565\(0) = '1' then
                \$1815\ := X"0000000" & X"7" & eclat_true;
                \$1814\ := X"0000000" & X"6" & work.Bool.land(""&\$1815\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1815\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1815\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1815\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1815\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1815\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1815\(0 to 31))) & eclat_false)));
                \$1813\ := X"0000000" & X"5" & work.Bool.land(""&\$1814\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1814\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1814\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1814\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1814\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1814\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1814\(0 to 31))) & eclat_false)));
                \$1812\ := X"0000000" & X"4" & work.Bool.land(""&\$1813\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1813\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1813\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1813\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1813\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1813\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1813\(0 to 31))) & eclat_false)));
                \$1811\ := X"0000000" & X"3" & work.Bool.land(""&\$1812\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1812\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1812\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1812\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1812\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1812\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1812\(0 to 31))) & eclat_false)));
                \$1810\ := X"0000000" & X"2" & work.Bool.land(""&\$1811\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1811\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1811\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1811\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1811\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1811\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1811\(0 to 31))) & eclat_false)));
                \$1809\ := X"0000000" & X"1" & work.Bool.land(""&\$1810\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1810\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1810\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1810\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1810\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1810\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1810\(0 to 31))) & eclat_false)));
                \$1808\ := X"0000000" & X"0" & work.Bool.land(""&\$1809\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1809\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1809\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1809\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1809\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1809\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1805_loop99401_arg\(32 to 63), \$1809\(0 to 31))) & eclat_false)));
                \$v559\ := work.Bool.land(""&\$1808\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1808\(0 to 31), X"0000000" & X"1"), \$1805_loop99401_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1808\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1808\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1808\(0 to 31),16),16)), \$1805_loop99401_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1805_loop99401_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1808\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1805_loop99401_arg\(32 to 63), \$1808\(0 to 31))) & eclat_false)));
                if \$v559\(0) = '1' then
                  \$v554\ := work.Int.eq(work.Int.add(\$1805_loop99401_arg\(32 to 63), X"0000000" & X"1"), \$1805_loop99401_arg\(96 to 127));
                  if \$v554\(0) = '1' then
                    \$1830\ := work.Print.print_string(clk,of_string("foo"));
                    \$1816_nb2\ := work.Int.add(\$1805_loop99401_arg\(384 to 415), X"0000000" & X"1");
                    \$1817_loop99398_id\ := "000000010001";
                    \$1817_loop99398_arg\ := \$1805_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1805_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1805_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1805_loop99401_arg\(32 to 63),32),16), \$1805_loop99401_arg\(64 to 95)) & \$1816_nb2\;
                    state_var598 := \$1817_LOOP99398\;
                  else
                    \$1816_nb2\ := \$1805_loop99401_arg\(384 to 415);
                    \$1817_loop99398_id\ := "000000010001";
                    \$1817_loop99398_arg\ := \$1805_loop99401_arg\(0 to 31) & 
                    work.Int.add(\$1805_loop99401_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1805_loop99401_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(\$1805_loop99401_arg\(32 to 63),32),16), \$1805_loop99401_arg\(64 to 95)) & \$1816_nb2\;
                    state_var598 := \$1817_LOOP99398\;
                  end if;
                else
                  \$1831_loop99399_id\ := "000000010010";
                  \$1831_loop99399_arg\ := \$1805_loop99401_arg\(0 to 31) & \$1805_loop99401_arg\(32 to 63) & 
                  work.Int.add(\$1805_loop99401_arg\(64 to 95), X"0000000" & X"1") & \$1805_loop99401_arg\(96 to 127) & \$1805_loop99401_arg\(128 to 383) & \$1805_loop99401_arg\(384 to 415);
                  state_var598 := \$1831_LOOP99399\;
                end if;
              else
                \$v564\ := work.Int.ge(\$1805_loop99401_arg\(32 to 63), \$1805_loop99401_arg\(0 to 31));
                if \$v564\(0) = '1' then
                  \$1844_loop99400_id\ := "000000010011";
                  \$1844_loop99400_arg\ := \$1805_loop99401_arg\(0 to 31) & 
                  work.Int.sub(\$1805_loop99401_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1805_loop99401_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1805_loop99401_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1805_loop99401_arg\(96 to 127) & \$1805_loop99401_arg\(128 to 383) & \$1805_loop99401_arg\(384 to 415);
                  state_var598 := \$1844_LOOP99400\;
                else
                  \$1805_loop99401_result\ := \$1805_loop99401_arg\(384 to 415);
                  \$1797_n\ := \$1805_loop99401_result\;
                  \$1798\ := work.Print.print_string(clk,of_string("rang "));
                  \$1799\ := work.Int.print(clk,\$1796\(1 to 32));
                  \$1800\ := work.Print.print_string(clk,of_string(": "));
                  \$1801\ := work.Int.print(clk,\$1797_n\);
                  \$1804\ := work.Print.print_newline(clk,eclat_unit);
                  \$1802\ := \$1797_n\;
                  \$v549\ := \$$1216_dst_lock\;
                  if \$v549\(0) = '1' then
                    state_var598 := Q_WAIT548;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1795_i\));
                    \$$1216_dst_write\ <= \$1802\; \$$1216_dst_write_request\ <= '1';
                    state_var598 := PAUSE_SET547;
                  end if;
                end if;
              end if;
            when \$1817_LOOP99398\ =>
              \$v553\ := work.Int.le(\$1817_loop99398_arg\(64 to 95), \$1817_loop99398_arg\(96 to 127));
              if \$v553\(0) = '1' then
                \$1827\ := X"0000000" & X"7" & eclat_true;
                \$1826\ := X"0000000" & X"6" & work.Bool.land(""&\$1827\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1827\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1827\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1827\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1827\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1827\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1827\(0 to 31))) & eclat_false)));
                \$1825\ := X"0000000" & X"5" & work.Bool.land(""&\$1826\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1826\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1826\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1826\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1826\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1826\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1826\(0 to 31))) & eclat_false)));
                \$1824\ := X"0000000" & X"4" & work.Bool.land(""&\$1825\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1825\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1825\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1825\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1825\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1825\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1825\(0 to 31))) & eclat_false)));
                \$1823\ := X"0000000" & X"3" & work.Bool.land(""&\$1824\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1824\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1824\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1824\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1824\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1824\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1824\(0 to 31))) & eclat_false)));
                \$1822\ := X"0000000" & X"2" & work.Bool.land(""&\$1823\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1823\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1823\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1823\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1823\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1823\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1823\(0 to 31))) & eclat_false)));
                \$1821\ := X"0000000" & X"1" & work.Bool.land(""&\$1822\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1822\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1822\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1822\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1822\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1822\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1822\(0 to 31))) & eclat_false)));
                \$1820\ := X"0000000" & X"0" & work.Bool.land(""&\$1821\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1821\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1821\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1821\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1821\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1821\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1817_loop99398_arg\(32 to 63), \$1821\(0 to 31))) & eclat_false)));
                \$v551\ := work.Bool.land(""&\$1820\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1820\(0 to 31), X"0000000" & X"1"), \$1817_loop99398_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1820\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1820\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1820\(0 to 31),16),16)), \$1817_loop99398_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1817_loop99398_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1820\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1817_loop99398_arg\(32 to 63), \$1820\(0 to 31))) & eclat_false)));
                if \$v551\(0) = '1' then
                  \$v550\ := work.Int.eq(work.Int.add(\$1817_loop99398_arg\(32 to 63), X"0000000" & X"1"), \$1817_loop99398_arg\(96 to 127));
                  if \$v550\(0) = '1' then
                    \$1829\ := work.Print.print_string(clk,of_string("foo"));
                    \$1828_nb2\ := work.Int.add(\$1817_loop99398_arg\(384 to 415), X"0000000" & X"1");
                    \$1817_loop99398_arg\ := \$1817_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1817_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1817_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1817_loop99398_arg\(32 to 63),32),16), \$1817_loop99398_arg\(64 to 95)) & \$1828_nb2\;
                    state_var598 := \$1817_LOOP99398\;
                  else
                    \$1828_nb2\ := \$1817_loop99398_arg\(384 to 415);
                    \$1817_loop99398_arg\ := \$1817_loop99398_arg\(0 to 31) & 
                    work.Int.add(\$1817_loop99398_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1817_loop99398_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(\$1817_loop99398_arg\(32 to 63),32),16), \$1817_loop99398_arg\(64 to 95)) & \$1828_nb2\;
                    state_var598 := \$1817_LOOP99398\;
                  end if;
                else
                  \$1817_loop99398_arg\ := \$1817_loop99398_arg\(0 to 31) & \$1817_loop99398_arg\(32 to 63) & 
                  work.Int.add(\$1817_loop99398_arg\(64 to 95), X"0000000" & X"1") & \$1817_loop99398_arg\(96 to 127) & \$1817_loop99398_arg\(128 to 383) & \$1817_loop99398_arg\(384 to 415);
                  state_var598 := \$1817_LOOP99398\;
                end if;
              else
                \$v552\ := work.Int.ge(\$1817_loop99398_arg\(32 to 63), \$1817_loop99398_arg\(0 to 31));
                if \$v552\(0) = '1' then
                  \$1817_loop99398_arg\ := \$1817_loop99398_arg\(0 to 31) & 
                  work.Int.sub(\$1817_loop99398_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1817_loop99398_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1817_loop99398_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1817_loop99398_arg\(96 to 127) & \$1817_loop99398_arg\(128 to 383) & \$1817_loop99398_arg\(384 to 415);
                  state_var598 := \$1817_LOOP99398\;
                else
                  \$1817_loop99398_result\ := \$1817_loop99398_arg\(384 to 415);
                  \$1805_loop99401_result\ := \$1817_loop99398_result\;
                  \$1797_n\ := \$1805_loop99401_result\;
                  \$1798\ := work.Print.print_string(clk,of_string("rang "));
                  \$1799\ := work.Int.print(clk,\$1796\(1 to 32));
                  \$1800\ := work.Print.print_string(clk,of_string(": "));
                  \$1801\ := work.Int.print(clk,\$1797_n\);
                  \$1804\ := work.Print.print_newline(clk,eclat_unit);
                  \$1802\ := \$1797_n\;
                  \$v549\ := \$$1216_dst_lock\;
                  if \$v549\(0) = '1' then
                    state_var598 := Q_WAIT548;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1795_i\));
                    \$$1216_dst_write\ <= \$1802\; \$$1216_dst_write_request\ <= '1';
                    state_var598 := PAUSE_SET547;
                  end if;
                end if;
              end if;
            when \$1831_LOOP99399\ =>
              \$v558\ := work.Int.le(\$1831_loop99399_arg\(64 to 95), \$1831_loop99399_arg\(96 to 127));
              if \$v558\(0) = '1' then
                \$1841\ := X"0000000" & X"7" & eclat_true;
                \$1840\ := X"0000000" & X"6" & work.Bool.land(""&\$1841\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1841\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1841\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1841\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1841\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1841\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1841\(0 to 31))) & eclat_false)));
                \$1839\ := X"0000000" & X"5" & work.Bool.land(""&\$1840\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1840\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1840\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1840\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1840\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1840\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1840\(0 to 31))) & eclat_false)));
                \$1838\ := X"0000000" & X"4" & work.Bool.land(""&\$1839\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1839\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1839\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1839\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1839\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1839\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1839\(0 to 31))) & eclat_false)));
                \$1837\ := X"0000000" & X"3" & work.Bool.land(""&\$1838\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1838\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1838\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1838\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1838\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1838\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1838\(0 to 31))) & eclat_false)));
                \$1836\ := X"0000000" & X"2" & work.Bool.land(""&\$1837\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1837\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1837\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1837\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1837\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1837\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1837\(0 to 31))) & eclat_false)));
                \$1835\ := X"0000000" & X"1" & work.Bool.land(""&\$1836\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1836\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1836\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1836\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1836\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1836\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1836\(0 to 31))) & eclat_false)));
                \$1834\ := X"0000000" & X"0" & work.Bool.land(""&\$1835\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1835\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1835\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1835\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1835\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1835\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1831_loop99399_arg\(32 to 63), \$1835\(0 to 31))) & eclat_false)));
                \$v556\ := work.Bool.land(""&\$1834\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1834\(0 to 31), X"0000000" & X"1"), \$1831_loop99399_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1834\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1834\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1834\(0 to 31),16),16)), \$1831_loop99399_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1831_loop99399_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1834\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1831_loop99399_arg\(32 to 63), \$1834\(0 to 31))) & eclat_false)));
                if \$v556\(0) = '1' then
                  \$v555\ := work.Int.eq(work.Int.add(\$1831_loop99399_arg\(32 to 63), X"0000000" & X"1"), \$1831_loop99399_arg\(96 to 127));
                  if \$v555\(0) = '1' then
                    \$1843\ := work.Print.print_string(clk,of_string("foo"));
                    \$1842_nb2\ := work.Int.add(\$1831_loop99399_arg\(384 to 415), X"0000000" & X"1");
                    \$1831_loop99399_arg\ := \$1831_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1831_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1831_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1831_loop99399_arg\(32 to 63),32),16), \$1831_loop99399_arg\(64 to 95)) & \$1842_nb2\;
                    state_var598 := \$1831_LOOP99399\;
                  else
                    \$1842_nb2\ := \$1831_loop99399_arg\(384 to 415);
                    \$1831_loop99399_arg\ := \$1831_loop99399_arg\(0 to 31) & 
                    work.Int.add(\$1831_loop99399_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1831_loop99399_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(\$1831_loop99399_arg\(32 to 63),32),16), \$1831_loop99399_arg\(64 to 95)) & \$1842_nb2\;
                    state_var598 := \$1831_LOOP99399\;
                  end if;
                else
                  \$1831_loop99399_arg\ := \$1831_loop99399_arg\(0 to 31) & \$1831_loop99399_arg\(32 to 63) & 
                  work.Int.add(\$1831_loop99399_arg\(64 to 95), X"0000000" & X"1") & \$1831_loop99399_arg\(96 to 127) & \$1831_loop99399_arg\(128 to 383) & \$1831_loop99399_arg\(384 to 415);
                  state_var598 := \$1831_LOOP99399\;
                end if;
              else
                \$v557\ := work.Int.ge(\$1831_loop99399_arg\(32 to 63), \$1831_loop99399_arg\(0 to 31));
                if \$v557\(0) = '1' then
                  \$1831_loop99399_arg\ := \$1831_loop99399_arg\(0 to 31) & 
                  work.Int.sub(\$1831_loop99399_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1831_loop99399_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1831_loop99399_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1831_loop99399_arg\(96 to 127) & \$1831_loop99399_arg\(128 to 383) & \$1831_loop99399_arg\(384 to 415);
                  state_var598 := \$1831_LOOP99399\;
                else
                  \$1831_loop99399_result\ := \$1831_loop99399_arg\(384 to 415);
                  \$1805_loop99401_result\ := \$1831_loop99399_result\;
                  \$1797_n\ := \$1805_loop99401_result\;
                  \$1798\ := work.Print.print_string(clk,of_string("rang "));
                  \$1799\ := work.Int.print(clk,\$1796\(1 to 32));
                  \$1800\ := work.Print.print_string(clk,of_string(": "));
                  \$1801\ := work.Int.print(clk,\$1797_n\);
                  \$1804\ := work.Print.print_newline(clk,eclat_unit);
                  \$1802\ := \$1797_n\;
                  \$v549\ := \$$1216_dst_lock\;
                  if \$v549\(0) = '1' then
                    state_var598 := Q_WAIT548;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1795_i\));
                    \$$1216_dst_write\ <= \$1802\; \$$1216_dst_write_request\ <= '1';
                    state_var598 := PAUSE_SET547;
                  end if;
                end if;
              end if;
            when \$1844_LOOP99400\ =>
              \$v563\ := work.Int.le(\$1844_loop99400_arg\(64 to 95), \$1844_loop99400_arg\(96 to 127));
              if \$v563\(0) = '1' then
                \$1854\ := X"0000000" & X"7" & eclat_true;
                \$1853\ := X"0000000" & X"6" & work.Bool.land(""&\$1854\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1854\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1854\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1854\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1854\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1854\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1854\(0 to 31))) & eclat_false)));
                \$1852\ := X"0000000" & X"5" & work.Bool.land(""&\$1853\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1853\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1853\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1853\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1853\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1853\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1853\(0 to 31))) & eclat_false)));
                \$1851\ := X"0000000" & X"4" & work.Bool.land(""&\$1852\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1852\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1852\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1852\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1852\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1852\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1852\(0 to 31))) & eclat_false)));
                \$1850\ := X"0000000" & X"3" & work.Bool.land(""&\$1851\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1851\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1851\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1851\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1851\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1851\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1851\(0 to 31))) & eclat_false)));
                \$1849\ := X"0000000" & X"2" & work.Bool.land(""&\$1850\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1850\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1850\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1850\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1850\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1850\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1850\(0 to 31))) & eclat_false)));
                \$1848\ := X"0000000" & X"1" & work.Bool.land(""&\$1849\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1849\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1849\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1849\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1849\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1849\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1849\(0 to 31))) & eclat_false)));
                \$1847\ := X"0000000" & X"0" & work.Bool.land(""&\$1848\(32), 
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Int.add(
                                                              \$1848\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                              eclat_if(
                                                              work.Int.neq(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1848\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.neq(
                                                              eclat_if(
                                                              work.Int.gt(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1848\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1848\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(64 to 95), 
                                                              work.Vect.nth(272, 32, 
                                                              \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1848\(0 to 31),16),16)))), 
                                                              work.Int.sub(
                                                              \$1844_loop99400_arg\(32 to 63), \$1848\(0 to 31))) & eclat_false)));
                \$v561\ := work.Bool.land(""&\$1847\(32), eclat_if(work.Int.gt(
                                                                   work.Int.add(
                                                                   \$1847\(0 to 31), X"0000000" & X"1"), \$1844_loop99400_arg\(32 to 63)) & eclat_true & 
                                                          eclat_if(work.Int.neq(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1847\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                          work.Int.neq(
                                                          eclat_if(work.Int.gt(
                                                                   work.Vect.nth(272, 32, 
                                                                   \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1847\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          work.Vect.nth(272, 32, 
                                                          \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1847\(0 to 31),16),16)), \$1844_loop99400_arg\(64 to 95)) & 
                                                          work.Int.sub(
                                                          \$1844_loop99400_arg\(64 to 95), 
                                                          work.Vect.nth(272, 32, 
                                                          \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1847\(0 to 31),16),16)))), 
                                                          work.Int.sub(
                                                          \$1844_loop99400_arg\(32 to 63), \$1847\(0 to 31))) & eclat_false)));
                if \$v561\(0) = '1' then
                  \$v560\ := work.Int.eq(work.Int.add(\$1844_loop99400_arg\(32 to 63), X"0000000" & X"1"), \$1844_loop99400_arg\(96 to 127));
                  if \$v560\(0) = '1' then
                    \$1856\ := work.Print.print_string(clk,of_string("foo"));
                    \$1855_nb2\ := work.Int.add(\$1844_loop99400_arg\(384 to 415), X"0000000" & X"1");
                    \$1844_loop99400_arg\ := \$1844_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1844_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1844_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1844_loop99400_arg\(32 to 63),32),16), \$1844_loop99400_arg\(64 to 95)) & \$1855_nb2\;
                    state_var598 := \$1844_LOOP99400\;
                  else
                    \$1855_nb2\ := \$1844_loop99400_arg\(384 to 415);
                    \$1844_loop99400_arg\ := \$1844_loop99400_arg\(0 to 31) & 
                    work.Int.add(\$1844_loop99400_arg\(32 to 63), X"0000000" & X"1") & X"0000000" & X"1" & \$1844_loop99400_arg\(96 to 127) & 
                    work.Vect.copy_with(304, 256, \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(\$1844_loop99400_arg\(32 to 63),32),16), \$1844_loop99400_arg\(64 to 95)) & \$1855_nb2\;
                    state_var598 := \$1844_LOOP99400\;
                  end if;
                else
                  \$1844_loop99400_arg\ := \$1844_loop99400_arg\(0 to 31) & \$1844_loop99400_arg\(32 to 63) & 
                  work.Int.add(\$1844_loop99400_arg\(64 to 95), X"0000000" & X"1") & \$1844_loop99400_arg\(96 to 127) & \$1844_loop99400_arg\(128 to 383) & \$1844_loop99400_arg\(384 to 415);
                  state_var598 := \$1844_LOOP99400\;
                end if;
              else
                \$v562\ := work.Int.ge(\$1844_loop99400_arg\(32 to 63), \$1844_loop99400_arg\(0 to 31));
                if \$v562\(0) = '1' then
                  \$1844_loop99400_arg\ := \$1844_loop99400_arg\(0 to 31) & 
                  work.Int.sub(\$1844_loop99400_arg\(32 to 63), X"0000000" & X"1") & 
                  work.Int.add(work.Vect.nth(272, 32, \$1844_loop99400_arg\(128 to 383), eclat_resize(eclat_resize(
                                                      work.Int.sub(\$1844_loop99400_arg\(32 to 63), X"0000000" & X"1"),16),16)), X"0000000" & X"1") & \$1844_loop99400_arg\(96 to 127) & \$1844_loop99400_arg\(128 to 383) & \$1844_loop99400_arg\(384 to 415);
                  state_var598 := \$1844_LOOP99400\;
                else
                  \$1844_loop99400_result\ := \$1844_loop99400_arg\(384 to 415);
                  \$1805_loop99401_result\ := \$1844_loop99400_result\;
                  \$1797_n\ := \$1805_loop99401_result\;
                  \$1798\ := work.Print.print_string(clk,of_string("rang "));
                  \$1799\ := work.Int.print(clk,\$1796\(1 to 32));
                  \$1800\ := work.Print.print_string(clk,of_string(": "));
                  \$1801\ := work.Int.print(clk,\$1797_n\);
                  \$1804\ := work.Print.print_newline(clk,eclat_unit);
                  \$1802\ := \$1797_n\;
                  \$v549\ := \$$1216_dst_lock\;
                  if \$v549\(0) = '1' then
                    state_var598 := Q_WAIT548;
                  else
                    acquire(\$$1216_dst_lock\);
                    \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1795_i\));
                    \$$1216_dst_write\ <= \$1802\; \$$1216_dst_write_request\ <= '1';
                    state_var598 := PAUSE_SET547;
                  end if;
                end if;
              end if;
            when PAR580 =>
              case state_var600 is
              when PAUSE_SET571 =>
                \$$1217_r_write_request\ <= '0';
                release(\$$1217_r_lock\);
                result568 := eclat_unit;
                rdy569 := eclat_true;
                state_var600 := IDLE570;
              when Q_WAIT572 =>
                \$v573\ := \$$1217_r_lock\;
                if \$v573\(0) = '1' then
                  state_var600 := Q_WAIT572;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1795_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var600 := PAUSE_SET571;
                end if;
              when IDLE570 =>
                
              end case;
              
              case state_var599 is
              when PAUSE_GET577 =>
                result574 := \$$1209_src_value\;
                release(\$$1209_src_lock\);
                rdy575 := eclat_true;
                state_var599 := IDLE576;
              when Q_WAIT578 =>
                \$v579\ := \$$1209_src_lock\;
                if \$v579\(0) = '1' then
                  state_var599 := Q_WAIT578;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1795_i\));
                  state_var599 := PAUSE_GET577;
                end if;
              when IDLE576 =>
                
              end case;
              
              \$v581\ := work.Bool.land(rdy569, rdy575);
              if \$v581\(0) = '1' then
                \$1796\ := result568 & result574;
                \$1805_loop99401_id\ := "000000010100";
                \$1805_loop99401_arg\ := X"0000000" & X"2" & X"0000000" & X"1" & X"0000000" & X"1" & eclat_resize(
                work.Vect.infos(256, 48, work.Vect.copy_with(304, 256, 
                                         eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1796\(1 to 32)))(0 to 15),32) & 
                work.Vect.copy_with(304, 256, eclat_vector_make(8,X"0000000" & X"1"), eclat_resize(X"0000000" & X"0",16), \$1796\(1 to 32)) & X"0000000" & X"0";
                state_var598 := \$1805_LOOP99401\;
              else
                state_var598 := PAR580;
              end if;
            when PAUSE_GET583 =>
              \$1795_i\ := \$$1217_r_value\;
              release(\$$1217_r_lock\);
              \$v582\ := work.Int.lt(\$1795_i\, std_logic_vector(to_unsigned(\$1209_src\'length,32)));
              if \$v582\(0) = '1' then
                rdy569 := eclat_false;
                \$v573\ := \$$1217_r_lock\;
                if \$v573\(0) = '1' then
                  state_var600 := Q_WAIT572;
                else
                  acquire(\$$1217_r_lock\);
                  \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= work.Int.add(
                                                                \$1795_i\, X"0000000" & X"1"); \$$1217_r_write_request\ <= '1';
                  state_var600 := PAUSE_SET571;
                end if;
                rdy575 := eclat_false;
                \$v579\ := \$$1209_src_lock\;
                if \$v579\(0) = '1' then
                  state_var599 := Q_WAIT578;
                else
                  acquire(\$$1209_src_lock\);
                  \$$1209_src_ptr\ <= to_integer(unsigned(\$1795_i\));
                  state_var599 := PAUSE_GET577;
                end if;
                state_var598 := PAR580;
              else
                \$1792_result\ := eclat_unit;
                result544 := \$1792_result\;
                rdy545 := eclat_true;
                state_var598 := IDLE546;
              end if;
            when PAUSE_SET547 =>
              \$$1216_dst_write_request\ <= '0';
              release(\$$1216_dst_lock\);
              \$1803\ := eclat_unit;
              \$1792_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
              state_var598 := \$1792\;
            when Q_WAIT548 =>
              \$v549\ := \$$1216_dst_lock\;
              if \$v549\(0) = '1' then
                state_var598 := Q_WAIT548;
              else
                acquire(\$$1216_dst_lock\);
                \$$1216_dst_ptr_write\ <= to_integer(unsigned(\$1795_i\));
                \$$1216_dst_write\ <= \$1802\; \$$1216_dst_write_request\ <= '1';
                state_var598 := PAUSE_SET547;
              end if;
            when Q_WAIT584 =>
              \$v585\ := \$$1217_r_lock\;
              if \$v585\(0) = '1' then
                state_var598 := Q_WAIT584;
              else
                acquire(\$$1217_r_lock\);
                \$$1217_r_ptr\ <= 0;
                state_var598 := PAUSE_GET583;
              end if;
            when IDLE546 =>
              
            end case;
            
            \$v587\ := work.Bool.land(rdy419, work.Bool.land(rdy461, 
                                                             work.Bool.land(
                                                             rdy503, rdy545)));
            if \$v587\(0) = '1' then
              \$1592\ := result418 & result460 & result502 & result544;
              \$1587\ := eclat_unit;
              \$1588_id\ := "000000000001";
              \$1588_arg\ := X"0000000" & X"0" & X"0000000" & X"0" & eclat_unit;
              state_var597 := \$1588\;
            else
              state_var597 := PAR586;
            end if;
          when PAUSE_GET410 =>
            \$1591_x\ := \$$1216_dst_value\;
            release(\$$1216_dst_lock\);
            \$1588_arg\ := work.Int.add(\$1591_x\, \$1588_arg\(0 to 31)) & 
            work.Int.add(\$1588_arg\(32 to 63), X"0000000" & X"1") & eclat_unit;
            state_var597 := \$1588\;
          when PAUSE_SET588 =>
            \$$1217_r_write_request\ <= '0';
            release(\$$1217_r_lock\);
            \$1586\ := eclat_unit;
            rdy419 := eclat_false;
            \$1593_i\ := X"0000000" & X"1";
            \$1594_id\ := "000000000110";
            \$1594_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
            state_var607 := \$1594\;
            rdy461 := eclat_false;
            \$1659_i\ := X"0000000" & X"2";
            \$1660_id\ := "000000001011";
            \$1660_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
            state_var604 := \$1660\;
            rdy503 := eclat_false;
            \$1725_i\ := X"0000000" & X"3";
            \$1726_id\ := "000000010000";
            \$1726_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
            state_var601 := \$1726\;
            rdy545 := eclat_false;
            \$1791_i\ := X"0000000" & X"4";
            \$1792_id\ := "000000010101";
            \$1792_arg\ := eclat_unit & eclat_unit & eclat_unit & eclat_unit;
            state_var598 := \$1792\;
            state_var597 := PAR586;
          when PAUSE_SET591 =>
            \$$1209_src_write_request\ <= '0';
            release(\$$1209_src_lock\);
            \$1860\ := eclat_unit;
            \$1857_arg\ := work.Int.add(\$1857_arg\(0 to 31), X"0000000" & X"1") & eclat_unit;
            state_var597 := \$1857\;
          when Q_WAIT411 =>
            \$v412\ := \$$1216_dst_lock\;
            if \$v412\(0) = '1' then
              state_var597 := Q_WAIT411;
            else
              acquire(\$$1216_dst_lock\);
              \$$1216_dst_ptr\ <= to_integer(unsigned(\$1588_arg\(32 to 63)));
              state_var597 := PAUSE_GET410;
            end if;
          when Q_WAIT589 =>
            \$v590\ := \$$1217_r_lock\;
            if \$v590\(0) = '1' then
              state_var597 := Q_WAIT589;
            else
              acquire(\$$1217_r_lock\);
              \$$1217_r_ptr_write\ <= 0;\$$1217_r_write\ <= X"0000000" & X"0"; \$$1217_r_write_request\ <= '1';
              state_var597 := PAUSE_SET588;
            end if;
          when Q_WAIT592 =>
            \$v593\ := \$$1209_src_lock\;
            if \$v593\(0) = '1' then
              state_var597 := Q_WAIT592;
            else
              acquire(\$$1209_src_lock\);
              \$$1209_src_ptr_write\ <= to_integer(unsigned(\$1857_arg\(0 to 31)));
              \$$1209_src_write\ <= work.Int.add(\$1857_arg\(0 to 31), X"0000000" & X"1"); \$$1209_src_write_request\ <= '1';
              state_var597 := PAUSE_SET591;
            end if;
          when IDLE409 =>
            rdy408 := eclat_false;
            \$1857_id\ := "000000010110";
            \$1857_arg\ := X"0000000" & X"0" & eclat_unit;
            state_var597 := \$1857\;
          end case;
          
          if rdy408(0) = '1' then
            
          else
            result407 := X"0000000" & X"0";
          end if;
          \$1578\ := result407 & rdy408;
          \$v406\ := ""&\$1578\(32);
          if \$v406\(0) = '1' then
            \$1582\ := work.Print.print_string(clk,of_string("cy:"));
            \$1583\ := work.Int.print(clk,\$1577_o\);
            \$1584\ := work.Print.print_string(clk,of_string("|number of solutions:"));
            \$1579\ := work.Int.print(clk,\$1578\(0 to 31));
            if \$v397\(0) = '1' then
              
            else
              \$v397\ := eclat_true;
              \$1581\ := eclat_false;
            end if;
            \$1581\ := eclat_if(\$1581\ & eclat_true & ""&\$1578\(32));
            \$1580_led\ := \$1581\;
            result403 := \$1580_led\ & "0"& X"0000000000000" & X"0";
            rdy404 := eclat_true;
            state := IDLE405;
          else
            \$1579\ := eclat_unit;
            if \$v397\(0) = '1' then
              
            else
              \$v397\ := eclat_true;
              \$1581\ := eclat_false;
            end if;
            \$1581\ := eclat_if(\$1581\ & eclat_true & ""&\$1578\(32));
            \$1580_led\ := \$1581\;
            result403 := \$1580_led\ & "0"& X"0000000000000" & X"0";
            rdy404 := eclat_true;
            state := IDLE405;
          end if;
        end if;
      end case;
      \state%next\ <= state;
      \state_var609%next\ <= state_var609;
      \state_var608%next\ <= state_var608;
      \state_var607%next\ <= state_var607;
      \state_var606%next\ <= state_var606;
      \state_var605%next\ <= state_var605;
      \state_var604%next\ <= state_var604;
      \state_var603%next\ <= state_var603;
      \state_var602%next\ <= state_var602;
      \state_var601%next\ <= state_var601;
      \state_var600%next\ <= state_var600;
      \state_var599%next\ <= state_var599;
      \state_var598%next\ <= state_var598;
      \state_var597%next\ <= state_var597;
      \rdy569%next\ <= rdy569;
      \$1737%next\ <= \$1737\;
      \$1646_loop99400_id%next\ <= \$1646_loop99400_id\;
      \$1685_loop99398_arg%next\ <= \$1685_loop99398_arg\;
      \$v511%next\ <= \$v511\;
      \$1664%next\ <= \$1664\;
      \$1744%next\ <= \$1744\;
      \$1682%next\ <= \$1682\;
      \$1762_nb2%next\ <= \$1762_nb2\;
      \$v596%next\ <= \$v596\;
      \$1577_o%next\ <= \$1577_o\;
      \$v447%next\ <= \$v447\;
      \$1666%next\ <= \$1666\;
      \$1834%next\ <= \$1834\;
      \$1683%next\ <= \$1683\;
      \$1633_loop99399_result%next\ <= \$1633_loop99399_result\;
      \$1637%next\ <= \$1637\;
      \$1646_loop99400_arg%next\ <= \$1646_loop99400_arg\;
      \$1803%next\ <= \$1803\;
      \$1797_n%next\ <= \$1797_n\;
      \$1698%next\ <= \$1698\;
      \$1735%next\ <= \$1735\;
      \$1730%next\ <= \$1730\;
      \$1685_loop99398_result%next\ <= \$1685_loop99398_result\;
      \$v561%next\ <= \$v561\;
      \$1756%next\ <= \$1756\;
      \$1765_loop99399_id%next\ <= \$1765_loop99399_id\;
      \$v579%next\ <= \$v579\;
      \$v557%next\ <= \$v557\;
      \$1719%next\ <= \$1719\;
      \$v413%next\ <= \$v413\;
      \$1811%next\ <= \$1811\;
      \$1703%next\ <= \$1703\;
      \$1821%next\ <= \$1821\;
      \$1640%next\ <= \$1640\;
      \$1633_loop99399_arg%next\ <= \$1633_loop99399_arg\;
      \$v553%next\ <= \$v553\;
      \$1645%next\ <= \$1645\;
      \$1627%next\ <= \$1627\;
      \$1613%next\ <= \$1613\;
      \$1712_loop99400_id%next\ <= \$1712_loop99400_id\;
      \$1578%next\ <= \$1578\;
      \$1707%next\ <= \$1707\;
      \$1814%next\ <= \$1814\;
      \result574%next\ <= result574;
      \$1755%next\ <= \$1755\;
      \$1677%next\ <= \$1677\;
      \result460%next\ <= result460;
      \$1638%next\ <= \$1638\;
      \$v512%next\ <= \$v512\;
      \result502%next\ <= result502;
      \$1815%next\ <= \$1815\;
      \$1771%next\ <= \$1771\;
      \$1684_nb2%next\ <= \$1684_nb2\;
      \$1660_id%next\ <= \$1660_id\;
      \$v550%next\ <= \$v550\;
      \result544%next\ <= result544;
      \$v507%next\ <= \$v507\;
      \$v406%next\ <= \$v406\;
      \$1844_loop99400_arg%next\ <= \$1844_loop99400_arg\;
      \$1816_nb2%next\ <= \$1816_nb2\;
      \$1791_i%next\ <= \$1791_i\;
      \$1843%next\ <= \$1843\;
      \$1817_loop99398_id%next\ <= \$1817_loop99398_id\;
      \result484%next\ <= result484;
      \$1628%next\ <= \$1628\;
      \result403%next\ <= result403;
      \$v513%next\ <= \$v513\;
      \$1639%next\ <= \$1639\;
      \$v540%next\ <= \$v540\;
      \$v517%next\ <= \$v517\;
      \$1665_n%next\ <= \$1665_n\;
      \$v543%next\ <= \$v543\;
      \rdy491%next\ <= rdy491;
      \rdy408%next\ <= rdy408;
      \$1597_i%next\ <= \$1597_i\;
      \$1860%next\ <= \$1860\;
      \$1852%next\ <= \$1852\;
      \$1787%next\ <= \$1787\;
      \$1705%next\ <= \$1705\;
      \$1593_i%next\ <= \$1593_i\;
      \$1853%next\ <= \$1853\;
      \$1831_loop99399_result%next\ <= \$1831_loop99399_result\;
      \$1765_loop99399_arg%next\ <= \$1765_loop99399_arg\;
      \$1710_nb2%next\ <= \$1710_nb2\;
      \$v581%next\ <= \$v581\;
      \$v427%next\ <= \$v427\;
      \$1732%next\ <= \$1732\;
      \$1585%next\ <= \$1585\;
      \$1736%next\ <= \$1736\;
      \$1594_id%next\ <= \$1594_id\;
      \$v471%next\ <= \$v471\;
      \$1678%next\ <= \$1678\;
      \$1592%next\ <= \$1592\;
      \$1726_id%next\ <= \$1726_id\;
      \$1697%next\ <= \$1697\;
      \$1594_result%next\ <= \$1594_result\;
      \$1850%next\ <= \$1850\;
      \$v425%next\ <= \$v425\;
      \$1603%next\ <= \$1603\;
      \$1681%next\ <= \$1681\;
      \$1725_i%next\ <= \$1725_i\;
      \result568%next\ <= result568;
      \$1672%next\ <= \$1672\;
      \$1790%next\ <= \$1790\;
      \$1782%next\ <= \$1782\;
      \$1649%next\ <= \$1649\;
      \$1623%next\ <= \$1623\;
      \$1856%next\ <= \$1856\;
      \$1825%next\ <= \$1825\;
      \$v539%next\ <= \$v539\;
      \$1622%next\ <= \$1622\;
      \$v497%next\ <= \$v497\;
      \$1583%next\ <= \$1583\;
      \$1792_id%next\ <= \$1792_id\;
      \$1751_loop99398_result%next\ <= \$1751_loop99398_result\;
      \$1751_loop99398_arg%next\ <= \$1751_loop99398_arg\;
      \$1611%next\ <= \$1611\;
      \$1734%next\ <= \$1734\;
      \$1724%next\ <= \$1724\;
      \$v469%next\ <= \$v469\;
      \$v470%next\ <= \$v470\;
      \$1669%next\ <= \$1669\;
      \$1835%next\ <= \$1835\;
      \$1693%next\ <= \$1693\;
      \$v395%next\ <= \$v395\;
      \$v431%next\ <= \$v431\;
      \$v559%next\ <= \$v559\;
      \$v433%next\ <= \$v433\;
      \$v495%next\ <= \$v495\;
      \$1673_loop99401_id%next\ <= \$1673_loop99401_id\;
      \$1691%next\ <= \$1691\;
      \$v481%next\ <= \$v481\;
      \$1716%next\ <= \$1716\;
      \$1601%next\ <= \$1601\;
      \$1702%next\ <= \$1702\;
      \$v432%next\ <= \$v432\;
      \$1625%next\ <= \$1625\;
      \$1857_id%next\ <= \$1857_id\;
      \$1745%next\ <= \$1745\;
      \$1685_loop99398_id%next\ <= \$1685_loop99398_id\;
      \$1848%next\ <= \$1848\;
      \$1830%next\ <= \$1830\;
      \$1742%next\ <= \$1742\;
      \result418%next\ <= result418;
      \$1692%next\ <= \$1692\;
      \$1581%next\ <= \$1581\;
      \$1591_x%next\ <= \$1591_x\;
      \$1776_nb2%next\ <= \$1776_nb2\;
      \$1676%next\ <= \$1676\;
      \$v590%next\ <= \$v590\;
      \$v478%next\ <= \$v478\;
      \$1670%next\ <= \$1670\;
      \$1739_loop99401_id%next\ <= \$1739_loop99401_id\;
      \$1653%next\ <= \$1653\;
      \$1699_loop99399_arg%next\ <= \$1699_loop99399_arg\;
      \$1587%next\ <= \$1587\;
      \$v516%next\ <= \$v516\;
      \$1837%next\ <= \$1837\;
      \$v428%next\ <= \$v428\;
      \$v473%next\ <= \$v473\;
      \$v467%next\ <= \$v467\;
      \$1712_loop99400_arg%next\ <= \$1712_loop99400_arg\;
      \$1607_loop99401_id%next\ <= \$1607_loop99401_id\;
      \$1715%next\ <= \$1715\;
      \$v466%next\ <= \$v466\;
      \$v562%next\ <= \$v562\;
      \$v501%next\ <= \$v501\;
      \$v593%next\ <= \$v593\;
      \$1659_i%next\ <= \$1659_i\;
      \$1827%next\ <= \$1827\;
      \$1617%next\ <= \$1617\;
      \$1750_nb2%next\ <= \$1750_nb2\;
      \$v435%next\ <= \$v435\;
      \$1851%next\ <= \$1851\;
      \$1743%next\ <= \$1743\;
      \$v573%next\ <= \$v573\;
      \$1788%next\ <= \$1788\;
      \rdy419%next\ <= rdy419;
      \$v520%next\ <= \$v520\;
      \$1854%next\ <= \$1854\;
      \$v565%next\ <= \$v565\;
      \$1805_loop99401_arg%next\ <= \$1805_loop99401_arg\;
      \$1781%next\ <= \$1781\;
      \rdy461%next\ <= rdy461;
      \rdy404%next\ <= rdy404;
      \result448%next\ <= result448;
      \$v429%next\ <= \$v429\;
      \$1694%next\ <= \$1694\;
      \$1840%next\ <= \$1840\;
      \$1775%next\ <= \$1775\;
      \$1629%next\ <= \$1629\;
      \$1712_loop99400_result%next\ <= \$1712_loop99400_result\;
      \$v480%next\ <= \$v480\;
      \rdy527%next\ <= rdy527;
      \$v509%next\ <= \$v509\;
      \rdy485%next\ <= rdy485;
      \$1778_loop99400_id%next\ <= \$1778_loop99400_id\;
      \$1588_id%next\ <= \$1588_id\;
      \$1841%next\ <= \$1841\;
      \$1817_loop99398_arg%next\ <= \$1817_loop99398_arg\;
      \$v459%next\ <= \$v459\;
      \$1792_result%next\ <= \$1792_result\;
      \$1768%next\ <= \$1768\;
      \$1632%next\ <= \$1632\;
      \$v521%next\ <= \$v521\;
      \$v476%next\ <= \$v476\;
      \$1598%next\ <= \$1598\;
      \$1657_nb2%next\ <= \$1657_nb2\;
      \$1644_nb2%next\ <= \$1644_nb2\;
      \$1696_nb2%next\ <= \$1696_nb2\;
      \$v438%next\ <= \$v438\;
      \$v555%next\ <= \$v555\;
      \$1718%next\ <= \$1718\;
      \$1796%next\ <= \$1796\;
      \$1844_loop99400_id%next\ <= \$1844_loop99400_id\;
      \$v424%next\ <= \$v424\;
      \$1584%next\ <= \$1584\;
      \$1855_nb2%next\ <= \$1855_nb2\;
      \$v456%next\ <= \$v456\;
      \$1619_loop99398_id%next\ <= \$1619_loop99398_id\;
      \$1817_loop99398_result%next\ <= \$1817_loop99398_result\;
      \$1642%next\ <= \$1642\;
      \$1619_loop99398_arg%next\ <= \$1619_loop99398_arg\;
      \$v426%next\ <= \$v426\;
      \$v397%next\ <= \$v397\;
      \$1689%next\ <= \$1689\;
      \$1847%next\ <= \$1847\;
      \$1679%next\ <= \$1679\;
      \result442%next\ <= result442;
      \$1844_loop99400_result%next\ <= \$1844_loop99400_result\;
      \$v537%next\ <= \$v537\;
      \$1783%next\ <= \$1783\;
      \$v489%next\ <= \$v489\;
      \$1809%next\ <= \$1809\;
      \$1849%next\ <= \$1849\;
      \$1607_loop99401_result%next\ <= \$1607_loop99401_result\;
      \$v436%next\ <= \$v436\;
      \$1826%next\ <= \$1826\;
      \$v472%next\ <= \$v472\;
      \$v434%next\ <= \$v434\;
      \$1602%next\ <= \$1602\;
      \$1792_arg%next\ <= \$1792_arg\;
      \result407%next\ <= result407;
      \$1778_loop99400_result%next\ <= \$1778_loop99400_result\;
      \$1761%next\ <= \$1761\;
      \$1708%next\ <= \$1708\;
      \$1599_n%next\ <= \$1599_n\;
      \$v479%next\ <= \$v479\;
      \$1748%next\ <= \$1748\;
      \$1800%next\ <= \$1800\;
      \$1823%next\ <= \$1823\;
      \$v554%next\ <= \$v554\;
      \$1726_result%next\ <= \$1726_result\;
      \$1626%next\ <= \$1626\;
      \$v552%next\ <= \$v552\;
      \$1824%next\ <= \$1824\;
      \$1695%next\ <= \$1695\;
      \$1699_loop99399_id%next\ <= \$1699_loop99399_id\;
      \$1739_loop99401_result%next\ <= \$1739_loop99401_result\;
      \$1747%next\ <= \$1747\;
      \$v498%next\ <= \$v498\;
      \$1650%next\ <= \$1650\;
      \$1624%next\ <= \$1624\;
      \$1839%next\ <= \$1839\;
      \$1651%next\ <= \$1651\;
      \$1667%next\ <= \$1667\;
      \$1673_loop99401_result%next\ <= \$1673_loop99401_result\;
      \$1652%next\ <= \$1652\;
      \$1646_loop99400_result%next\ <= \$1646_loop99400_result\;
      \$1802%next\ <= \$1802\;
      \$1777%next\ <= \$1777\;
      \$1671%next\ <= \$1671\;
      \$1757%next\ <= \$1757\;
      \$v453%next\ <= \$v453\;
      \$1720%next\ <= \$1720\;
      \$v563%next\ <= \$v563\;
      \$1749%next\ <= \$1749\;
      \$v549%next\ <= \$v549\;
      \$v585%next\ <= \$v585\;
      \$v423%next\ <= \$v423\;
      \$1805_loop99401_id%next\ <= \$1805_loop99401_id\;
      \$1699_loop99399_result%next\ <= \$1699_loop99399_result\;
      \$1842_nb2%next\ <= \$1842_nb2\;
      \$1774%next\ <= \$1774\;
      \$1723_nb2%next\ <= \$1723_nb2\;
      \$1633_loop99399_id%next\ <= \$1633_loop99399_id\;
      \$1612%next\ <= \$1612\;
      \$1829%next\ <= \$1829\;
      \$1785%next\ <= \$1785\;
      \$1733%next\ <= \$1733\;
      \$1773%next\ <= \$1773\;
      \$v515%next\ <= \$v515\;
      \$v439%next\ <= \$v439\;
      \$v551%next\ <= \$v551\;
      \$1688%next\ <= \$1688\;
      \$1582%next\ <= \$1582\;
      \$v430%next\ <= \$v430\;
      \rdy545%next\ <= rdy545;
      \$1822%next\ <= \$1822\;
      \$1654%next\ <= \$1654\;
      \$1786%next\ <= \$1786\;
      \$1828_nb2%next\ <= \$1828_nb2\;
      \$1798%next\ <= \$1798\;
      \$1778_loop99400_arg%next\ <= \$1778_loop99400_arg\;
      \$1857_result%next\ <= \$1857_result\;
      \$1660_arg%next\ <= \$1660_arg\;
      \$1641%next\ <= \$1641\;
      \$1769%next\ <= \$1769\;
      \rdy449%next\ <= rdy449;
      \$1857_arg%next\ <= \$1857_arg\;
      \$1726_arg%next\ <= \$1726_arg\;
      \$1610%next\ <= \$1610\;
      \$1804%next\ <= \$1804\;
      \$1754%next\ <= \$1754\;
      \$1759%next\ <= \$1759\;
      \$v465%next\ <= \$v465\;
      \$v531%next\ <= \$v531\;
      \$v508%next\ <= \$v508\;
      \$1643%next\ <= \$1643\;
      \result490%next\ <= result490;
      \$v564%next\ <= \$v564\;
      \$1656%next\ <= \$1656\;
      \$v437%next\ <= \$v437\;
      \$1586%next\ <= \$1586\;
      \$1760%next\ <= \$1760\;
      \$1813%next\ <= \$1813\;
      \$1721%next\ <= \$1721\;
      \$1680%next\ <= \$1680\;
      \$v522%next\ <= \$v522\;
      \$1668%next\ <= \$1668\;
      \$1831_loop99399_id%next\ <= \$1831_loop99399_id\;
      \result526%next\ <= result526;
      \$1746%next\ <= \$1746\;
      \$v560%next\ <= \$v560\;
      \rdy443%next\ <= rdy443;
      \$v475%next\ <= \$v475\;
      \$1588_result%next\ <= \$1588_result\;
      \$v477%next\ <= \$v477\;
      \$1607_loop99401_arg%next\ <= \$1607_loop99401_arg\;
      \$1631%next\ <= \$1631\;
      \$v582%next\ <= \$v582\;
      \$v514%next\ <= \$v514\;
      \$1772%next\ <= \$1772\;
      \$1739_loop99401_arg%next\ <= \$1739_loop99401_arg\;
      \$v455%next\ <= \$v455\;
      \$1580_led%next\ <= \$1580_led\;
      \$v587%next\ <= \$v587\;
      \$1605%next\ <= \$1605\;
      \$1820%next\ <= \$1820\;
      \$v468%next\ <= \$v468\;
      \rdy575%next\ <= rdy575;
      \$1801%next\ <= \$1801\;
      \$1660_result%next\ <= \$1660_result\;
      \$v556%next\ <= \$v556\;
      \$1861%next\ <= \$1861\;
      \$1764%next\ <= \$1764\;
      \$1836%next\ <= \$1836\;
      \$1838%next\ <= \$1838\;
      \$v558%next\ <= \$v558\;
      \$1738%next\ <= \$1738\;
      \$1630_nb2%next\ <= \$1630_nb2\;
      \$1579%next\ <= \$1579\;
      \$1805_loop99401_result%next\ <= \$1805_loop99401_result\;
      \$1729_i%next\ <= \$1729_i\;
      \$1751_loop99398_id%next\ <= \$1751_loop99398_id\;
      \$1722%next\ <= \$1722\;
      \$1618_nb2%next\ <= \$1618_nb2\;
      \$1795_i%next\ <= \$1795_i\;
      \$1758%next\ <= \$1758\;
      \$1658%next\ <= \$1658\;
      \$v519%next\ <= \$v519\;
      \$1784%next\ <= \$1784\;
      \$1763%next\ <= \$1763\;
      \$1588_arg%next\ <= \$1588_arg\;
      \$1616%next\ <= \$1616\;
      \$1808%next\ <= \$1808\;
      \result532%next\ <= result532;
      \$1655%next\ <= \$1655\;
      \$v594%next\ <= \$v594\;
      \rdy533%next\ <= rdy533;
      \$1765_loop99399_result%next\ <= \$1765_loop99399_result\;
      \$v523%next\ <= \$v523\;
      \$1604%next\ <= \$1604\;
      \$1711%next\ <= \$1711\;
      \$1663_i%next\ <= \$1663_i\;
      \$1636%next\ <= \$1636\;
      \$1799%next\ <= \$1799\;
      \$1810%next\ <= \$1810\;
      \$1831_loop99399_arg%next\ <= \$1831_loop99399_arg\;
      \$1731_n%next\ <= \$1731_n\;
      \$v474%next\ <= \$v474\;
      \$v510%next\ <= \$v510\;
      \$1594_arg%next\ <= \$1594_arg\;
      \$1615%next\ <= \$1615\;
      \$v518%next\ <= \$v518\;
      \$1717%next\ <= \$1717\;
      \$1706%next\ <= \$1706\;
      \$1606%next\ <= \$1606\;
      \$1789_nb2%next\ <= \$1789_nb2\;
      \$1600%next\ <= \$1600\;
      \$1770%next\ <= \$1770\;
      \$1709%next\ <= \$1709\;
      \$1673_loop99401_arg%next\ <= \$1673_loop99401_arg\;
      \$1704%next\ <= \$1704\;
      \$1690%next\ <= \$1690\;
      \$1619_loop99398_result%next\ <= \$1619_loop99398_result\;
      \rdy503%next\ <= rdy503;
      \$1812%next\ <= \$1812\;
      \$1614%next\ <= \$1614\;
      \$v412%next\ <= \$v412\;
      \$$1209_src_lock%next\ <= \$$1209_src_lock\;
      \$$1216_dst_lock%next\ <= \$$1216_dst_lock\;
      \$$1217_r_lock%next\ <= \$$1217_r_lock\;
      
      
      result <= result403;
      end process;
  end architecture;
